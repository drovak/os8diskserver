����   � *?>22
%? 
      <
>!"52	=<(*"<;:2. 2">(/987	6988	*,.   548#38: '2++'2+: +#;$'2/9+'2/9: +#.5  >(/                                                                                                                                                                                                �+&@ٔ�MA    ���                                                  ��7��@� ���Ѝ��� t�W��?���� ?V������������� 2�K���Z֩A�?�����s�
��� �v���? ���?�� ���� ���� �������(?�~�!�c(�����(?�~��c����6������&�,� �
�&����!b��  ܳ�*�b��f!�,�   ھ�+�b��Ӛ!�,�  Ղ��}�������}/�����l��  �(?��?���������|)�ظ � ҁ�������� �f����Ɗ��/�ۨ���(��!�����J���H/�(����Ϩ,�"F�ۀ��F�,
.
���h���
��&,� F��ۀ��"�b�j���-���/Ȁ�� � .�b�j�9�J� ��|��{����,�$ۭ�t�c�%\�� �AP�CrR� Ђ�� H���  b� ����+�&��r-�h--r.-d�-���z�..7 
.
�z---t-�"���O�*���� ���T� �����&��� ���/f�ʈ/�(�"�����J zD/./��8�K � ,,b��/�,���K堮��c��@��b���� /��@�v��?�?`������ ׀��  !�����&��&��l��
     ��~!����(?���6�6�6��ˁ"¨���&�	&�&F>�	7�J� ��&�&�&���b�n�˚t��ˀ��٨�����t������٨� ��/���Jٿ�D. b ��l�Ub!�l!t��/�����!� �������! |	���(���H/�� ,,b� ��{����,�"(���@.��/�,��@.��/�,���K':"ȇ�q�9�/���{z$�8��)�7��6)q��5&����9�/����)�) &�)�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3 �
����?  �W����