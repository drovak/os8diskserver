����    �@7$> .: 
./
 ./41!  8>(*+?7<: 7:8 
0>(*);7<: 7>? .:
../
-./
?  
7"9
8"9.1
  0&0!*;: .9  0+ 0>0&0!+=<(/<;<(/:9<(?87.?  ?7>(/65/U5 ? 24>>                                                                                                                                                                                                  �@ٔ�MA�':�!�  X�ŀ���    �     � �� ���  � @  �� @�    I�     � �     k   ��� �   �^�UB��� R@� � ����dB� ��(�?��s�@: ��M��8m�e��a��$���g2�� ��`���f��?��������@�JA�J���!B��&(?�B������6��c!C�7C�J�6��/@����"�j��)��)�����������F���������iÀ��ꒊ����/���/��"c(��������0F����0��&�0�&�*  x�/?��� y?u�1�9� ��S�_jQl�l��~	 �Q���  	��A���� �Oj��jd v�O"�p
�
��� H  �y |���D�PQU��A	 S � ��D                                 �����-��ڠ����r��r���������������������� �  � ����������ʈ��������J� ���-������נ/�Ѥ�����? a� � �͍�߃���� �����Ju &�+��w��n 6��+�(��+d_2(���(/������� ��
&
(?�(�`�z�����b(bi(l�4�lv	�?�������2�ހ���? ������� N�������� �H/��O�������j8�   ���ƌ�+	������!����̯�&�����"��hˍ���&��&�톖����ގ���"��* ���O� ��F.���+��   	���F�H��	�������j �
'�	a� �����᠎��&��(���������္���� ������	��F
�������h�� ֚�������������yz'z{'��݃�݃������-��݄��߉�g��-��ݎ���������J�j�o��V�0�-�+�+D��,��(߈&�0!.10&�+�('J ��+�t�c%� �)����ɥ��%� }�9���N��ߎ��ڨߑ���ߓ����+��B���a������-��� �⨩�����������⯭����P� �(��(����  &!̻��� �����&!����(���(/���(���� � ���-�����'�t���( L"�|���� ���g{�������j �)|����?r �����8                                                                                                                                                                                                 