��� L C    �B �?��b�r�TU�(�!�r�b(���J!:���k�8�   � ��_9��� ^�{7����4E)��ʉp�4E)��ʉ'��a�������E9�ρ �0E)� ˉ ��&�&�	&(?���	T9/(�¢�1bB��+�/�5�5b5c��5Ks c�J
�4H.>�                                                                                                                                                                                                �������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ  �
��D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �      �8���}���v	P�nݏ_��F� ��&8H.�����H/C�/�ڮ�/����"�i���&�!.��/�Ȩ���}Ɉ  ��b�bW�ԉl�@�|"����"��o�'����"����J��b(���}Ɉ � ���k��hB�?�D����Ի �?�"���V�"�����'�N��PTB 0��� ����� � �,�` VV�!�۠/�F����۶��r��x|&���(��m�/����(��m�(��@��|&��y�����m(/��������z�� �"�b� �F.��+�(/���H��bV���������m� ����⨉�� �۠/��� 8f��0(���O頮�)�����? 8����W�f'2��pD�F�&�`>E��� E��
���	&u&A�.��&��r��/ @��f�����|�&�J��|�&O������ݨ*���C 	�u�C !��H��	�r� ��F�?����r��	�'|�� /����"��s��{   �(?��B6� � ��$�֚��pWgJ��(���o p�x�݈����/���}�� %����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� �������  @��      8bD8��&m F���@/�ԦP���J�כ��"��O���������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�޴�����2X��(?�
�

��������ς����o��R1��D��� N E��D� �@C劀���	��T P�ل�MA	O���� 0���/a�   ���f�	&�	��J�g�v��KV�e�� �@� �? ����]���aOY����&7�B!!⠌�!�6]Z9Xc��c'���b��&��7��b��/����naa7�!.�`bc�t��!&`!>S"���O0�����b!a�@��a�xM>]]s��/�O�MT�a'�!.cc7]rG�* a�`b�f�?��`!>&�2��d��          � � ����6��6���H  �� >u������c{�J�����t��7��C?�F�0�F'��0��c_���t�6�>0bJ�8�c{(����m"�m�m�&�m"�d��&�l鈐  0���k �&�9 O��J���`/���������n��&� �    Vx��DW�b��o��P��Dd#pD 8��/�8�������m�(��@��|&8&8J.8����(���H/�J�V�8&��,� � ���'�J>
��H.��J
��������u��(��!�瘨Ϩ�H��{ J
�?H.��J
�������r��{8��8�c8V�k      �G�w x� g�P�@ ��� ��\�_"VU�2d                                                                                                                                                띓��@��������Ӎ� ������?�!�}] c�� @ ��U�