���  @  B 	/   	    	 	    (	) 	 	 	       ,    	     	   	 	   	                                                                                                                                                                                                 �����&��&ތJ���  �#&���(�����������������������(�����������������(����������������)��)��)!�  �"� 0���'��)��'��)�	�$b&%b'�b��{ � �_ ����dB��F V�f�fE�v �尭U��U�P��U �@�����)��	�b�i����'�!%⠙�'�/�����)��[������������'�!�&�&$�&�"`���������(� �bJ
�
����&��"�!i   �
" �  `����&�"�bJ
�!��b�l!>�Á�ϙ��J�����)�����[�WW �	p����1gR�E�"g̴U� U �f��[��'��)��������3�6�)��)��9��)��9��)�(?�����)�(?�����)!.�(?�����)��
�O���r��d��J~�)�Ê��&��B��ry�/4@�~����� �=kR��b��b�@n�u�N�*u��� �M�/|��� ���y����O��g��w��w�og��e��U��e �f�fR�E ��F�Á�� ��F�2��h ������������� �666�<�� �
�'���  ��!�"  �	�<br�!�
�<���� �             ��h�ֈ��)�̋ b

�
���)��H���&�P.��/�󩀀�������G���f����@���F � &�&(?��7��������c(��c�z��K��b��c(����b�$6%�b�&!>��&.�%b!$�$�b��c����/��"�n�&%6�?�%�������	�h�J��"c(���J.
���d���� �       Nfabfcdfeff$%  �
n')�H��T��� �f��l	 `          �
�             �
�#ǁ#Ė&�!�ʀ�� �� �� ��� ���(��(� ��b�bcf"H��F����"���������� ��
>

�ױ�ױ�� ��(���(����(׫�� �� �� ��(�a�c�� �khPoH��� �?� ����� ��PAA�H�H�A3:XS%V������1��^ � So�#R�� @T��TXV`��dN�� �(�3ɇSL�h�D�ԃT�ȟ � PF0��L�`�PR0S�#P��5 N 	ϋ���8�R� AN(�8�`�8I� (�A)3L�`R�$�%�8(M`�E3Ճ��7T��D��  �D�ԃT�����HLS!Ճ�8��1� E�����HLS!Ճ�8��4τV�C_! �5ND!	ϋ����4 ��)b�����J����#6�#+��B��z��(�2����"d!)b�\�[�&������@�� ���t���v`�v��U