���CD �E � ��$8$  !=-Z$l8 a  &&2&2	') '$(%/>>/!>?8 {"/*[8?>/=;    {*8�B E:54), }-	 <=���������                                                                                                                                                                                                                                                             ��������É��l��� ��ͨ��É� �������|؋<�&6���� �  �������� �,��������ɀ ���	��� ���?���J����i� �� ���hӀ��!��� ���ͫ   ��É���.����� ��$� � 8��8�kH_T���J0 ��j�we(9χ�������2�����̼�� 7�����2(����/�����~��x�q���"��s�/��"��{����ɀ ��� ������'��'������Ÿ��y���(����(� ���n큜_��K���Ŵ��������'遼��s���"ʉ|�^�( �� ���d��- ? ����dw���q~N�R��RYy8��Y�6�/�J.��(����&��É�������b����B�j��/��6�&��)wwt(?��C�z�� ����������9� ?��(?�ɶ� ���   (����6۝ �����)� ��g���&��B��   ����d� � �� ������7Yy_��  �`�o< ��
Ҧ� � T	� �h�n �	�� ` �   n � @Ć �z�� `T������ �
� � � Ė �k责o    � � ��o ��� X ��o  ��N�Ħ �k � ����� ���� `T�� T	�訤o  ��NƦ T	� ����� �w ������ T	� 訣o  ��NĆ ��訣o�@  ����� �� � �   � � �Ć� � ,� 谤o   �<�訤o  ��N   � �? @(? 0 ? @ H 	ĥo  @K�� . 8	� `Wm�          ��<���� ��<���;����L���� ����U��U��U��U��U��U��U��U��U��U��U��U��Ufff!$f+2f5<f?BfEHfKRfU `   � �   � @   �     
G 
A(7 (
G 
�       � �G�#G   �     
G��A(7� �G�G�G�#G27�-      
G�A(7��G�G�b�b�Ѿ    ���� ����� ��N� ��t�� ��}� ����� �°N� ��£� �A�>� ����� ��>� ���L���� � @��� ���d·6��K � ���!.�b�b������9� ���&��6�����������&������ Ap��������MNU j�Y�=ЛR�� �	�	ߨ/��2�i�ߒ����2����ߒ�����8�(�(�(�*�٘��8ߨ/�F>ȕ��ݠ/�����bgww���(/��(���(/��(���/���������7�����K�'� �G� ������N�/���� -�p�����/�	%��!��k#Y <�����0͎� �� ���"��f��i�O� ���"`��/����D.̯bH�����$����"����b�����+       �����/�բ�bb�b��c��������&���    	�β�{�	  ��6��ǉ�����s��{������� nֶM����T�{�<���	�������	�� f�b�n��f���(���/���" ��(����/���暀����"����H.&/���t���������&� ��"����?���h�����h̀���h�����)���6��6��C麚 �	b�ڛ�����빀� � �=蛮��S����?�	���A�]�� ��/����/��b�c(��(��������︻����6��&��9   �
C٤�@����F����������D� �   !�(?�����D��� ���?��?�˻��� ���� �(����i� ��ߛ�c�/?�ߛ�&� �   �^�]T  �p���� �N�]�x �&�(���p.oN�� .�{ �@�����P.�/��K���
 ��&�&t��� ��(/���(���(/����Ǹ�����(���(� ����<�����&�����F���|�"(���k ���{���#� �-��pߧ�W� �`��� կ
F� ���6�������/� �� �b

�
���(� ��(�������� �����������(�(� ���i���������/��������/�в��(����/���!��&����̯k ���4�l�<����<��@����/�ԋ    �����ꋀ��!����}] ]��� ? �M��+���������6��)� �����)�������cb�����)�)�)��� �	#�� �	+�� �	3��r:��:P�: �4 �T��G �J F��: �
   � p!����N��NJ p ��l�׊��(?����������� ��2 ���J��+      �` �� T*pL�K ��� ��d Z �	�� � ��/� ��ŀ�  ������ �	� �� ��6��'��)�&� ���4(����� ��b ����É�� .�/��� ���(���(/�����ǉ����  �����i����� �  �������  루��  ������  �	 � �	  ��D�p�������  ��W�ͳ� � ��G��"����� �	�����  �	�Ԁ��	�� �� �� ��  (����/�ؾ���(����������  �   ��6��C�b�����2������    ���	��b���k�R� �������ҋ ��|���ỉ��w���+����8����� � ����?��p�T*�#; �Z  ��l�?���&�'�|����{ ��lC�(Ϧ��(����/����ǉ�˒�K �����i(����/����y����r�i���(���cǂl��� �����b�b�l�9J
�d�9F���逞�D��   ��M�ǀ����#�O ��]g0͎���@����D� ���  � (���(/���@�����'�����®�n&����� ���b ��߁l��<��/�ɤ��B��� � �B��� �� �!���@n��"�����)� ā ����� � ���r��y�c�n&��'���6��'� �����ÉJ�
����+�H/ �.���+ � Y� ǩ �� �� ��6��N�6��C��d����d�/��?t���� ���˛��E�����<���O����:�� ������7��������&��2������� ��
>����&۠?���
     �̲��r���۴�(����Ͽ���<��~��r��r��r�G������������� kyP�]��T� �(����bF�����b��&��É����)��b��,�ޖ�J.����b���݁l���JP�����P��"��&��"��c���@������"ہlۉ<àn� ����B��� ������)���Z�������@�         � /��
�   ��߀� K�NjZT�]��f�hg��F���� ���?�������FN���&��,��|��C����������i�����i��������(���� �    ��� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d������ ����� ���� � (����B���ǉ�� ��������9��s������C���z�� ���ɀ 5���K ���� 5����� ���s!� ���)��)��� F�� ��É ���@� ����f������{����?���d��� ��L�����ѝ� `   �ʌF��:�?߇( �TN�<0��?  ��/�����b��b��g�'Ӝ'�����y�&�|���xD��r�   ��c��������Ө?��0�����0��s(����tĠ?���������� ���N �	���(�����<H����)��+ ��bg�J������|؞� �-�����N0 ?� 8G ���Џ���k��ߗ��                                                                                                                                                                                                �Xct�c � �����,c�t@���� ��L�pl��@>Eo3���t@@ҐFt@	%%�aRc) D�t��0l 	�3C �	���� 9A�2P N� 4n -�K ���e;SWn �� E�pJus �խHt�c�%\�� �AP�CrR� 8�)  �    �
��G���b��h�����'�������� �
����i� T�������  �������̀@ � ���d��2����ӊ����P.��/�٨�!���0��O�٨����J�ъ���ǀ�������   ��J�
>

�堮��c��@��b���� /��@�v��?�?`��؇��� � ���F.����&��� �挀'8� ��/�����t����F.��+,0�58�;=�@C�GL�PÚ�#R@��A�T A� BP� A3@�b� 0�# U �� �MA���5����5BR1 �BR  y� dgi�kn�ru��E��D�O3�5S �QS RU��A@�(D�T2� 0���   (���(/���������Łl����d�(?�����b�����!��Ȼ��>����F.����0��'��0(���H.���!>��<��������� ����� � ���b��$@����&���(���F.���+    ���{ �����ƪ��A@�0�:��o�&�)#�:�8����P� <� �Œ��	8��0MN0 ��3��R`N` O�5�NB�PTB 0� 5��T ��4:Q ��4��CE:1 ��4�	D�0��0��EO3� @` �� 5N��M�@�hN� �PN�M��`6	I3 �UL`!��CN�!�          S	PRQ�	A� 0CN���MM��BT��USB	�#S�� ��ϋ���8��4� @��GLN� V�σN�`�a�4ԃՃ� 0Ń��C XQS %�N��TR���O����C �VC`� 0���H��C �DLN!M`�8��CA�	�	��RC! �Q 0�̓A�3N�`�R�� 0�D�M�����GL*���O�D��N�� 0�D�Ʌ R�	5� 0�̓A�3σ΃������C��N�!XCL �8�U �# LP�5 � @�D�̀Ʌ R��3 �DC��0O�#�D�V�C@!�΃DPC%�H�U�$��;-���-�̀F� DT  �� �� @�  � PP��@̓0� 48C � P	��	  @B�DRD0 �  5�@P 0� E � ��@��@�DσD� �$ 0��@ � P �   0# A�L	�3 � ��  ��  � Ҡ �� �� �� �� �� �� �� �� Ȯ �� �� �� �� �� č �  � �� S U @d AP�3�8 �� ��&(?������������ �꒢��b�b��x��(����b��/��������"�������j���� ���(��(� ���G��"���� ����  ��ŤؓD���&����͎������� �
��� ���d�(?ܹ���J ����	 SրD^]}����`�� ��"���E��                                                                                                                                                                                                