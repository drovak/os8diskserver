���� �   H�  &-	  39>6/6v 
"> -9 	>*<*9 
&>*
%*9 
'>*
$*9 
#>-;-  7                         3;98= 1> 1.1 %.>4v? 6   6 4                                                                                                                                                                                                                   � �m   S      �� �                         �          � �s��
         *     ? @� ��   �?����� ��`��00U=�� �$_��U��U��d��̍��][�T�d��E��v����dC�z�u!�q ��������������������¤���;�&S�#�����4�H �4C F���@�� 3b��� �"��h� �����`���� �O��ҡ�� �
 � 1%`�K� "ƾ&@�龀1E�i?�� �4A   bD � "��� �&� !����r�ny�ϒ��r	�b
�b �l	�<
 t�n��j���X�2��/�$�&%f� �sE0s�{4< (���&�%	!�P�KM�����P��4r@J�M'Kl�������Ȩ����"D�S	sJ>���� �                            ���6IA.Wo�:A.V9�(/� �YX�9 D��98"�N��Y�9!.:K{� P�lt�6u�6w�6� �   ���NH�4�k9 0��'��� P	�k   3�/�4��F	&�		c�	c"b`"�N�(	c(���b`�␓�Q)@�'n((&'D.)(b"�@'�))&(�"(&@)�	&(�F���&4@ J
����n�a	�! K�  �O��ҡ��
�4@ J
����Pn�ݑ߀�1E�i?a� �(Siv)6r�/�(�)�|s�0�s'� �� ���'���� �  �H �⨂� �'��N��&��"����&�H�HH"�������   ����(/q�� ����j��/�����������"���!�˖&<��䖙"�����&��K��K�� �� �� �� �� �  ��Á����	�&�&Ӥ�45&P6�K�4�k:�0M'�'_��r�r�r�r�k�����0��@4< ��&��+b�3 �Bhz�3C�0e963;:3`K� � b�?�C&�#�l ?�|# '�O �J��� Z	%�/����L�%�/�[����}%B���;0&�/&.�[���i��1f"#f�1�11c�(/⎢(���B���"�J.�/�#����A�*#�/�"����,1'�#������O�i�)P���1KZ��\Z�L�[K�Z��\Z�L�[K�ǒ	�+�P?� �x� xc���� �w y��2x �����x � ��4&���H��� � �!���� �"c��i@ JN9 �& �"�OiR�6TK;Y�? YZ[3\�33(o3O����OE����3zA���� �� �� �� �� �� �� �� O����c�,��oA Tn��� @�&�D��%H/N�%$b��$G"(��@N�$%bH$䢍�%�+ �	�x�utsvss�sj���o �4�A  D. "
�c
:6
6
86��`.
�?�8�!A�HA�"bQ:�:n(F.�b��c:96�,�4��FP.��� L!�{>@K��g� L	?JK���L$�$�"�N�$r&$�"csGb�b	�b
	c
��JK��rs �M�������%�(����/���X%�Kk �3_i9"�K�@���9�/�I�AW�o��"�hYia���9�JOKY�@F�����%Kk�J�F����9�JK �"H.f:C��d=�"bH����Q"��+ :��;�&��1�K�9r�K�:A.W�(��X �!�I�Vp�YX���b��/N9��K�H� J

���b=���sJ>P�sK{ 1(Gb'"b"�(/�@�1.('d�"��� w�N�� �`.�/Nϔ�<��3Kk  77B!���N� 7'�>�T.�Kk� P,J)�J){�{�  s�0����� %�`�� �\j��q���(/KX�9Ib
�i
9t�K�ɯG9An:V)b+�-(/������98"���+X)9�JN,�+b�)e9!.:K{��b(K�!{���/kI�AW�o�9Yi  bF�/>?" J)9�JK���� hK��/���J���b�b{cH?稯K��k�K��hK��J)��JK�p�_���Ƞ���Kkr�/���K�� = 2�e��/�2�d2��=02�'��/������;�& ���l���D�
 �� ���k    �Ġ/�ţd=�2�b ��2�,�ųŭJ��b;�&��* �� �ľk    r���Bt#!v�(����D���ƴ�1�iƛ ��� � ii�� U)�ݛ�v�v rF�  b� �F��f��{� C �iAU���c �	N�sJ>���NK��v��� �	vsSJ��N�K� S	v�6r�/��Á�� i	���(�?�++b��/c��f�vv7�C��hCJ
�J
�f�{h���g � j�$��%��&�KӹK�� h	Nr�����-"�T�gj� ��r����+�&���I
&9&�/K:����;�&v:c�
�9OK9��K�h��g��� j$�U%�U&�U����)11C��/���1r{�2�k�1-2���1�81�J��(�K{oU_� �  b��/�h�N{�r�/�g�j � e�� R)�� s������u�X�����u�x!>u`>y�?����cy�`z�c�y�[� @��T� s����T�ꈸ tvss�s�� ]	j�+ ]	}$"���%�/�_��%����`�"'fX#�$!.#bX#�'.'d�%�#%&' &"b���]z��}�%"&_"�����<��z�`��\<�� �    ]q�]t�%�&4�i\ǐ�%�(�������/������]w����w%"���\w�%�&�]�w\)w�)<]yw%"���\t��q�]t��_�K����w�O�����\t���?K��<K{\<�K���N�\q����w�)KP����?
{ %(K�Ȣ�� $�aK� ���f���"%b(���`�$H/�$o$ N������
�()f�%"%%b(&����(�H(�).)�i)�"a&�(��#n(�"a%��� ����J "�%#b&)bD���(b����n�"d���%�b&�k  �/ � � ��p��˂����j�����<�z`���<�]}��]�z�)������z�)���z�)���}�(� ������ ��� �O��@
�  ]}��$��ai�}�� �%�/�`���� �Р/`˛ �	����]}����������}])z\)}$$ ��z�)<�y�$"$�k � �                   �	]}��<�%�/�\�<�y}])}.�\i}�)]z��&��#�� ��z������z������}���/�����C�K �%h/�F�($�!�(&���$&f%�k$�&$]i}�))]�z\)}�))�z])}�)]z��2��/��z��,��}��5�]z��$&a�z�)8��� ��
�O ����H� p�w���6�_�t�H�p�U�����,~
LD`�n���o�k9r��䷊�l��� ��` `�xR�  P�vq �U �  @ �����/�� �$`/ǀ��آ(��@��$@n%H/�%$d�%�$�k�� 0$%&&�b$^i� ��"6�Q)��sH%�$n&!f^K��;@���Ȟ�# ��O���$� ���v.�/��0�b/�l��'%(/����ީ�$r����ϚߕJ�]�m$�Z%�&.b���!0�@ ��H/���Ʋj�ϚưJ�m��$�!���ř�'&.�/�ߦ��*:/� $����Ϛ ����jh��p�z>�_���� �Ҁ�] ��
��"@���/"!��0(/ ��@����j��)��J����ߒ@��!��0�/������� >�0b ��訾O�懶�!0�`���.⠶��ŀ'�/����(�n�'bH!�&%f@��&�(�(&%�$��-�/�不��� !�%b(&b)�i������"�i����i�.��J������������ �/o���� ��{ ���� �   �/� ���O�䨪�
�������� �� ~��l*$f&�`%�fҚ�*�D�Ϛ]}�\̚^ʙ}�*ɡZ��D�����dà��+bƨ/Ұ�#F.#D.ͨ*#�$!!��a.Hq� ������d��� �
�]�m �;���һ 
�      P #�+��(/������h+�"@���o��KF �b*����+�"����`�U��  �������_� m	��9��ɀ�+]U� m	��9&)&"&6$a.'$&'%b"(b%"b(�l��'��'�*��(��ֻ �	���#(b����#�)D.)(b(�!%b����#� '�]�f��"a.%/�@�%�i!@/�@�&O�%&b&�$ N%�*%�k���$�(&�%�i&a.&o ��-  �t�	Cb��b�	���J��˚  s>2s�{ m	��9$$&�"f%�/$�h()&�"�&�b%%b��!��#D���� �$$&���/ ��'&) /�!��)�)���@"�&"&%��.�"b"�!�'�J�)�"/�@�&.")b���a�&n�D� m	��9!$�$(ba(��&�!�b��jҀ&� �%("����"&�%�%�%("%��&�&�"�J�]�(����� m	��9�(¨��%�/�$�a'�`��!��'�$�h���������   (b��(.()b)�"�' N �J� �!D.!&b&�%.%�k   %b��%.%&b&�!�$ N �J���� �mϓ��π&���	DA�0��  &a.&n%a.%�k )a)�(�a(�� �@"�!!&)�&&&(�%%&�a��� ""'6�"�  �(�h")6� �%(/&(/!�/�ڮ% /�&�����ܪ!�k/ �m���'�$)b&(b%�d��� m	��6$�'�%���x&�'��L� ���K�������l��� "�Ȳ�!�%@n(%"��% n!!&�%��b�p$�$�i�$��è�A3� 0�$�瀻NN�_K�N �sJ>�h�Kk�K*������D k��Rt�vfyH���,���?,++bR�+�"���+�"(����/�+�eg�� � ��kr������v!>t�?���Ri����f��vv7�ܠsE0?s'�s�E>s�zkВ��&+e)tv7f��4�� �4J.
<�� �7�"�N�7 6�7�7 b�վ����xMK{�$��%��&�Kɴ sH����K�� D�"�K�`.B�/�<���`�␒���*`.��/�����`��K�;&K �w 4   #               s�0F�`��������N��Ѐ Ѐ �                                                                                          