����  � ��	           		  ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                    �+&@ٔ�MA � ���L �    F  �  �                        �0�    �
�	�   �
� ��   �Ī��A � � � Z
    �d@�@�@@I@@�@�/@  ��� ������������  ��K� ��� �� �� ��                         ���< �<�<����<i$τ��01f�2&��&��&�*&�+&�,&��&��/�2��*s+0t��/�2��*s,1t,�D+�D�O�2�*@N�.�@n�.�@n�1����0�/�����b� n( n��t��J�&<7�<B�-)�EHv� �      �   ��� u (��|u |)�ظ� ����h��xp h   ���93i5��8:�6�-K�-/˝����խ�<�J0�D=i���93i5��8:�6�-K�-Ӥ���ٜ<�S0�D=i��� 	���� 9A�2P N� 4n -�K ���e;SWn �� E�pJus �խHt�c�%\�� �AP�CrR�	1G                         )���95i�8:6��K��/����Ԏ�Ճ�<\�0D&=���9&5��8:�6�-K�-Ӣ��5��8�E'K�-/˝����խ�<�e0�D=i���9:i6�-L�-M�-���/ԝ����<�n0�D=i���95i�8:6��N�����խ�њ<w�0D&=� � ��b���� /��@� �P? ?`��؇ ޱ������95i�8:6��O��/����Ԏ�Ճ�<��0D&=���9&:6�FFb�L��M���ݣխ5��8F��N���ݠ��/ҝ����խ�<��0�D=i���93i5��8:�6�-N�-/˝����խ�<��0�D=i���9Lb�:�6�-P�-���/ԝ����<��0�D=i뀲!�l!t=��!�z�<"�i;)eO"7"���93i5�� :	6F&F�-K�-ӎ��Q��/�ӈ�Մ�<��0D&=���9&35�� p:6�FFb�K���ݫխF�-R�-Ӳ��F��S��P����T�/�/�ӈ��UШ��ա�<��0D&=Λ 2�&wաڅ���4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� �Ș"���93i5���:�6F&F�-K�-�VҠ���F��R����W��խ5���F��N����V�/�/����Ӫ�Մ�<��0D&=���9&35��p~:6��K�������/ɝ����խ�<��0�D=iπ��- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0I.3���93i[�&[�&\�&B�&��&5��8:�6F&F�-K�-Ә��5��8F�-K�-Ӣ�Ԥ�ƚJ�^�`_�_^�__�^_�ǰJ_^�_Ȕ�_�^_�ɺJ_^�_ʔ���� �       �����ݢ�!|�ԫ�����d��6� �   �ۢ�݂��d͊���  ��� ���d�� �v �J
�
��(��H��ĳ���9�b��b
3i:6�Ffia�����9:i6F&^f�a������1��e������ �� �� ��  <	�
�A<��0�D=i� ��@�Uu��٨�@�Uw��٨� ���6��Iy�O�Xi �����  y\i d	a	r�� ��ٛW+,wX ����� �@e�`	 b�a	 r�Uy��R�����@L@@F��D�<��.�)b�c�g&d����94i5��8;�c�-K�-/˝����խ�<�J1�D=i���94i5��8;�c�-K�-Ӱ���٨<�S1�D=i���9;icF&F�-���M�-����5��8F�-N�-ɠ��/�҈����ս�<��1D&=���9&;c��L��M�����/�Ԉ����<n�1D&=�� aYr���D� K��D���95i�8;c��N���݋խ���<w�1D&=���9&g�&45�� p;c��K�������/ɝ����խ�<��1�D=i�����<ڜ.)�bc&��bgdk ��e���@�r�+ ���d��6�WIX ����� �  \ �c��e�c �d�^ �d�` �]r�� ��!l��{�/�{��&,���   ���7-� �                                                                                                                                                                                                 ���=��C��Ԁ ���6��C��d�E#GHf��E�G�JH�BG n ���G�(����* I� J�Jb��h   �C�Hb�rGvHEg� � @C�cּd��6��B��jC.CCb�/C�n�.��dȼ�    � ���/�ʣ(��@����/����ʤ��J���&�/���'�/�ʤ��6� � �`b�� ��խ�8&0!.��b�6b��j ��խ�8&1!.��b�cb�8c��-Ԟ�̲Р����-Ӧ�Ԩ��8Ա�J��� �    (���80b ��884ԴK�L�(9k (���81b ��884��K�L�(9k   �8&0!.�<i>8�A��A8���J� ��8&1!.�<i>8�A��A8���J堰 ����Rxp@   �EKr�/�ɠ�ӈ�Ԋ�Հ� &!��"�Ύ ����Db!D�?@f>9�A)�?& @�>9�A)D�J����k Y&!̳"��X�&!̹"���렮 � ���f�Bb��b�o�@n��"�����?���?�J�(/���������@�/徢���A����D�@�?�k�,���� �    � n������ 5	�8F�-K�-ӈ�Ԋ�Հ� Z�F��M���ݕԭ�խ� �5��8F��N���ݣԭ�խ� �5��8F��N��/����Դ�թ� 5	�8F�-N�-���ո��<���ˆ  ���	�d	�6�
.

��؂�Ί   �(���H����* ������ ����*�&,!��"���?����� �k�]O"�62�u艅EN��O�	5E�4��wAN2�8D�C#A޷ ��C���E߀G��t�07���;�`NCP��#RTO�#��w��	�S� p N�T  0 �`  �  ��X`�0 Q`6 �T`!�TE�  ��TR`�R   � �΃��CP�  ������Z� �D%נ3  ��TR`	� H  � �H(��0� @�H`�0 Q`6 ���%��� 0�TR`O�   � R��F E` �X�R1S` ! `N� T�`` �     �  � އu�ݐ`  �  �ް| ��` (  � އN �8MN"߀�� �DM�P��HG1L*�����D