����C� C<(+.5=282	$/842/ e4 ?=?>?%   ? ?8 >6<���������                                                                                                                                                                                                                                                                                                                         ��b��b��b��f�(?����&��&(?�������k��R����(�!.��/�����/������ ��� � ́��φ������ ��7��B�����t�O�͈�5�� ��(?�P���"�����"��b��&�Ɉ�� ���"��b��b��k�J��� ���	�O� �0��Mօo�L��2c����� �7�
���`�������&�!>�i�|��0�c�b����(?�!.b�c�� ��&��������� �f��&C����'�"�br�& ��c�!>�?�������������1( P �0� �B�2�O�p� ������w����?��b�f�&�è�����&�/���b��&�&�)�(/���(���!.�l�)�¨��͙J�b&��#���� ����D����J�"H����� ����!.c������� �&'!>&�Z���J��&� �C�{��?P���I�� � ��0�c�@������8����Ȁ��/��"�i�����a.����&���ŦJ�&������"����)�J�Ê!.����������� ��>������h��0���� �����b�bD���b����)�J� ����崁�!����;����& gK�pI�]������"&6������������������F� �� ���ј���!.�������� ��&������ ��[�6��r܉�����)����	@n	�2�����i�6� ��ޘ�	��	�9���� �� ��(���,ޚ�f]��̿�̂B� Kw�XX;��?��o��   A.����/���F�
��۴	�	
&�D�ܲ�������� �!.����!.���ט������)�+ / ����	�"	`O�(�� ��&	!.�b �d!.
�b��b	�k ��
�� � ���+I��4N (L���2- �      ��������������@�X�KBx �(���c�����i�/��
���(��d�������0J
��(��&�������)�ĸ���)���Ę��/�D���&��� �
����� D���� ����!>�bվf��b(��@����d����� O���ߢ� ������OsEm; �X���;
��M� ]�� ��"b	�b�	�
b�*&�?����� ���q����׉����ਭ���(q>�8���hq>�8D�J
$��	d���� �����?�����!�67'D�J� �b&"�k �ffb	c&	6�"�i	�?���&� �M�_.	  &!����� ������b�����������
ɀ(� ���{ �!Κ�?�������(��(��(����K  �扱ø�h �� �!������ ��)�)� �D����?���� �

�
�� ���"�c�(�����J��B��{��3��C҃T� E� r	<? ]���@ ހ 碟RCč � ���; ����; j�*�S�UCm2 ��N  a�SmS ]�G1L? ]G1L* Mt~ h REq���Y��MA ֆE�tO�#]UL��	5�8D  �D R�C� @]��8�	E�8L@!]��8�4�8L@!]��8A	�8RC!�T VC`S�8V``	��@�@6�8XNR �D �N �B]R0]]Y0�N%�L%]G�PA��0��3C ��a.������ ��&�8�c�a�� /����c�a�0� �(������c�!�/��"�,� ��(��"(���(/���H����,ݛ��"��k@  @���� ? F �������֮��������P�����(?��'�&��)�(/�������J�&�&�)�/�֮ /�/B�����������"����b��c(��������*��iT ��̢��r�b��c��� ��آ������������,���������� ��O�����I���	���1����