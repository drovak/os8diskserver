����  �. . 00000000  .	  ; 	8: 18	 *%
.
/%
3
4%
;
<%% 1	
%%%# 0000   0000  : 0000   : 0000%#.  00000000  .  9: 18%                                                                                                                                                                                                �i� �;`.:" � ���/          �   ��?; ?G �8� @�??�p    d   �3 ��  � �� �� �� �� �� �� ˨ ө  ������ !       L��!��  D� � �    �)�"�X!x��
<��  � x肁�^� Zx�,D� ���

c��b

�
�菐(� � � (���@/������ ����*� /������&!̥���"�
�?�������  � �6� ���
�$0�c#��"0�c��J.��
���&��H�'�.����&��H�']�&��K      0�� �bD�.Hs�b �J��"�*n &��,�m�����.&.�&�-��+'/' 0f��ގ � ���&"b!⨤��*��(�6&3&"��(?�&�!�ʬ����.# ��1'b(" �&��1�-I����%11�-! ���&�?��-LM��?��-LM��?��-LN�M��?2�L�MW���� .��c�LKrJ p�a��0�!2�z�!.�/���"gk�� ���1D[�1f[ �&	&OD. �OOb	t��� �1�-��� ����� ���Ԩ�����ڡ�ݲ���R���S&�Р�����U����� .فlJ 0�(��R�Tٚ! �s�g"�n�bQF�u�7� �P(/i �Oy��m�L#� ٔC �bbb	bcQ	cPQb!P⠕��J������S�b������b� c��V��_�a�!��"����0ƿ��e���e��He�f��.�&�-� ,a._,,̻ �S.�1�T�S* QYiTopY)QtuY)RxyY)1��Y)S��X)c�`00 �`00���00�cB��H�00�00� �K  �S���1.TSb*RYT���"YR���"YQ���"YP���"Y1���"YS���"Xc�`P00� �`00�� 1�0�0 ȁ �0�0c�B� 0�00�0 �� �D.�1�T�YT���"Yb���"Xc�CP�0,0 �R���D�0�0 ��X�cL�.	8��; Xc�NQ�	��;  0�1c!!bL��9��&!�J�F.(��  �
(�,� �0�iw> ��㙂��h�6����b����/��㨠��D������>�*�!&�!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0�H>                                                                                                                                                                                                