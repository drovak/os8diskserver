����  � 
/ ?<0 ? 
=3?  5?, (?=> ==   * 0'4	 8 :"���������                                                                                                                                                                                                                                                                                               ��@v&xş��C ���G �� �                                 6 0����))K ��~��}����7|�01�7�@ �� �� g�1Iv @�!߈� ��?���� ����
s� �� �(�/�}�  (� �BA0�����Q�!� ���&{ɀ{)��(b!'�{֒�'�(��&{��z �b!#�{��z��$#b@ �$�/���y)by!��/�{��"x{��"!%�wb%H/��%@/��v!.b%b!�{��z �!ba.$/�%�!.%$�!�%&ut'st�"&)��#" ���r�a.$�/�� z	 q�J
��{���*$&���}��-}� �(/��&$�%�t�"bb%pk)�r�b�}�on) ��&�����bb%�hp �"b&� ���m�(l����k�jig0 &� i��-jg�(�
u�&&!�/�}�js��
h%2!��&�&!> ?������J{�gk��n}֚ ��-)f�k"H��n����e��0��{�ze�e �ƽd�ec"(���bB(l�a@.`/��D.DD�&_"ｈc /�{��"� ����� ^&.�] _����« �\[)�6�ZB[�(��YJ

���X@�ۊ W@Y�V[)� �!��&��� ����UF_�[z���� ! f�T��S��)�RQ"�PbO�~�N��� !.H���N��� h��ݟ�����|����J �"�dn)���M�  /�%�!h�"O'��=����@��|��}������N���h�?��T�� ����e�����U�' /Lh�!(�(&DK�TJ���@����k�&e�-�����J� ��O����{��gћ�P`�p�`  �� �P��2X�`6ԠL`
 �� 3���%Ѓ`j�L ` ��C���C��NTR# ��DX��C�����  ��T�TT?(X=E��1HN�� �����  PX� 5 - NτT�D��@��2 � 0�TR`R��D��NTR# ����#�5��� 0!&�(�({i�"�(c('(!>%�/�)�d *�x)&�J�T�   I�-�h�HO'�����߱G���ݫe��hӝ|�S"��� p ���v&xϐ�	HA�1�� 7|>�������	w�k�x�ԃՃ� 0 �8�8�8����D7)8)���|ly���a�S��*���{�x9��E�� �                                                                                                                                                                                                