����    �3# /  82# /  2> 2!'2/ ; 	#9	8	0, ; 	#9	8	0,   !<2/9  &5��������������������������������������������������������������������������������                                                                                                                                                                                                              
 @ٔ�MA�� ���L � /BNX � �v  �wqp� � �������������         �7��x       �    ��<          PX�iq�@�/��z�g �����? ( W�(�X��Z֩A�?����s�
��� �v���? ���?���R��` �P������/��� ��������ɀ�� ����� �� ��x����
���F.��b
�Ⲳb��������⸳{o���K���뼁���'��'����ˁl��'�&�&����]����ښ ��h{

������ u (��|u |)�ظ� �� �(?�r�� ,
�����6�������6��B (�
�

� �般���)����� ����K ���)��   �� ��
��b

�
鯪��?���� �?� «��
.��´�)»�ՠ�)�δ���  �צ��&  ��,&���d�� F"��!���H�� �JH� �/J�� J            ���
.	�!.	 /�		b!
�!.b	
" /�
	" /
�	" /�
"	 /�!⨸�
&
&�*�&�	&�
&
'
	�٢�r�{ �!�	&�&��!� �	�J������ ��7����6����ۤ�� �/2��y2K.)��2���� p�6��7�� ��� (� ���b���������.�!�⨜������3 ��ܒ<"c��b����&���@/�â@���J��2�;�����������������D��
� �
�/���>>!.�/�>�D���>>b�?&Ł�����-�%2`n/�@x�r������an�%͘dC4f�b�??@	��E��� 0�H>�(C!&㠀�#�?�����(/�"'2� 0`&%7ڐ$$s��/�$���/���))�2ȡ�ސ#y�@**s�!�(/�����-�/����+&�	&*�0�����&��
�
� ���
� ���
'	�J���?����8 � � ��� � ��� ���d�� �v �J
�
��(��H�� �-/ (����� ��*7*����6�+�	i��H	��J����2�v@�����d� & n�� s! �&�@ ��%� �奈����n�x%��d�- n%��p� ���N����| �/2��y8���{;�d��':&(;&il��j��:�!8� ��;!.9�/�l��m�����R���\L���3��3�3(!>&�?�����(/�"'2� 0P(!>%�?�'���������(��"2{��D8'���(!>%�?��A(���(��ר =�3��@�5琠�� '�H��=O�'�;���'����$'7�(�((s W���;�'(?�ݦ3 ��@�5琠��'"w;@�4��@�5;� (�!&���3��@��4��@5�;���=�8(c!&㠊��$�����������)�63 ��@����8=D� �=�n��}��)�6��"!Hﹴ�ȹ�4 � @�����D ����r��i���)�6�8�88b�2���b]�/��!�=&F.�&8>&9?&�_���Xr�k��R  �ߴ��
{�/�{��&,���   ���7-���U \����O��5����/�'�8�F ��2����{�:R�!��/�����i���)�6�8�H��8�j�<䯮�I3y�@5�)�4i �@�J�� � *b���U)&)�J*�J�˺�/��I�/g˛zb�I"�/�����t��sw�=!.q��T��� ��X&�IРb����@ � "b���"7� 8������'�!$㨩�)�63 ��@��'��;K�'�R�) �P'�!$���)�64 ��@��'��3� �@��͠���&'W((S Wਲ��#�@#��%����"';Y��4� �@���@� IЀ���&O��Ϣ"w25� ��2���{\f��O�3��@5�)��3i �@Ԛ���� p �� ����,�-�ny�k���������"������p0n0�J//b,��ި���(/�΢���/-"-/b,,&���k�/� ,�,/b -�-�h����,�/�ި�'��Ps��I���� �!�������)�������޻ ����%��$�����2��2����?%	%%� ��?  ? 3����ҝ�֮0�-��݋֮0�-���נ�L�Ɲ�"�y��2��2�0�-���2̽ר����n"	&	t���"2{��?�':� �/2 �y�2{.)Ȳ{IV~0�-�խ����L�Ɲ�"w2 ��2־0�-���2־0�-���נ�L����"2{o�}20�����2���Ш��"(w'2{񀀮�̀!>��� ��À�0*#>�-��&�9֠��=�:ր�M���2ˡNy6@/�V�������6‭���0*#>M >�-ŭ�!�� N��=��B�c��M�9��:�������ΧN6�@��V�����N6�+���ӭI���K���o ����������� � ���� �� @�@2Iv@���� G����*�
��� ��*@2*�{�� �.Xn//b,��/�H.䖟�./BH/�/�  ������,�������!�ﳪ.H.
�0.b�&�	&�
&	
t³��ؠ��f�H.�� ���H.�����+�    ܠ�y2K.)�!K9):��6)7���(��'9ܻ      ���7� ���6�+ ��2���\����'I� ��2������� ��2��������� �!%����o��x%��d����o��� �x%��d��!� o�?��Ǻ�&?�&��&��&��')!>	�b
�n+&�<Py	�J�&�R�'�9 P��(Q0R�) PǛ
�J���            ���?���b��b��n��4�n)!>	Sb�Tr�v8(/�!�'�R�)! �P9����N(Q0R�)! �P9����U�
�n�U�
�n+&��!P��?�	���
�J�\��!>S�/�βO ��2�����T�' ����M� ����s!S����'j�8�k��]�-�����-~՛@<�� ����ƙ����!�!%в���!�! �!2	��������J �����t�'��K �
��c��c��d���P����M���� �      ?�&?�& �P��R�� ��Py� � �-/ ����*�����)�Ų�ƽ~���@��խ�����-~ڛ �/@<� �瀮�-����̭���������խ�@�J��H?��8�������'!>$�?�'�(XX"8v;@������^ǔ�*�0��/�)��3i �@�i�=�;��)�64 ��@����=�j����b	)c!
�?�&�ð	
�JP��Ā�'!>$�?�'������ BC�D��Ћ EF�G��؋ �� 6����l���D�(C.B, ��G�(F.E,  ���&��� �	                                                                                                                                                                                                