��� Cm �D2 v "���������                                                                                                                                                                                                                                                                                                                                                                          ����B�l��&�� ����ہl��D���������@.�/�ozN

���&���� �  `����"��b�D��  ���&��&����������Д�c�J
��

��J��0��d��0�(/���� @�������c(���� �0 ��Z
�d�6F��K����f��P�S� ��&��&����(���  ����� ����y��L�����������خ���� ���l��?��(����&�F.�����bP�Ⱗ���̍ �   ����K ���?���������������ȟ��"����(/��튁�9� ȋLȨ�  �9?P@��;PU� �:�P� �!�淸b��k � ��l��&��/����O����F.�බ7�J.
�����r��d��J��)��������d��'�O� �   � �   ���ŉl��0��&�?� ��,��/�˃�� ��/�ǲ�����г��&��+��]�T	���@ a�/�	�a⠀� ��}����� K ��� ��������������9� �� ���&�'�&�&�'�j �	�/��������c��c@�����z
�
���i���    �		��&ض����������&�à����������X.����r���'�����n&��������PGU�`+fD]�D M��
T:���g���'�y�&(?����Ԣ��������?������  ��0�����)����'��0�����0�����0����>�����?��� �������?����������)�ߙ��i�ȿ��ԄJ   ���� �    ����9m	���`�Pǥ� ��� W����������� �Ԁgi�G��&�v���� �(/���(���&�"@������&���f��fрo'�B��/��������'��B����'��������'��)���&�'�J������'��)������c�/ߠ�&���z   �������`�������� �� U�l�r�\e�OM� ��&����&�(?���  ��I   �	���&�J� ��F���
@�ဠJ���&��&��9  ����r����[����� ���'��f���n�s�����"����'w��y�w�r�7����� �	� �  ���@  �  �  �  ���� 1y �4�J�'����;u���       P�@�����  P     � ��               n �                                  ������&(?���a��o���J�#��{ ����أ���������/BD���������K�J��� ��l��G�Y������ �ȟ����/��t������c(���� �
���� �
��2����>����f����� ����b� ��d�	6��Bc	t���]�S�`X��6R�RC�HS� A &���!��� ����/���������/�ݫT������L��4Ȁ�퀏���t;� �	������&�������;P�s�``�`C�RQ��C � N  a�SmS ]�G1L? ]G1L* Mt~ h REq���Y��MA ֆE�tO�#]UL��	5�8D  �D R�C� @]��8�	E�8L@!]��8�4�8L@!]��8A	�8RC!�T g	����;��	�������͚(��Ơ/����Ƣ(���&� �(/����(����������Ƃ������ �@������&��)�J����~��

���c`��(���h��Ź���������� ��)�ٚb�������H�����v�T.� ����	��\ m��IWg�8;���`����g ��&
>

����� ��(���������H.� ��(/��(��(��(�H���"�����"��k@������� �� ?���ʂl�	� ���� ���i
�   �������������  �   
��$�-9�IX�gt��b�B �       � ����  �����V��?@ ��3��C҃T� E� N`!�S�3	����]q��CL�TN�� 0RC�H��C � N�	���3TUL�@VC_�8R�C�HVC@�AC�T����� ���7]#GLN�R`N$,XL_! � DRC!�T�����]�#TX��C ���7Z �^���w��w��������c(���� ���J��������&�'�6�����  0����  �������r�뙠����{ �(��!� ���0�&�?��� �Ӂ,��r��rߋ|� ��a>�?����S��O�����������C���_�B�އ��f�D���?;��]d�K�����G��&������� �����6�	&	(?���&�	�b(��`��/���~��7!.�/�/��!�b!�b!��"�����S����2������grwr�u��(����렞�&�	�����`H]�ՃR� ��+ ���9Ҁ��:��۔�����u��݄����r(/�������s���ؙ����H�����x���
  ��&��� �� Ж������������)��/������� �	���,��r��w��� �m�#]��	8�8-�O�sNI%� 0��3��C	��-�O��N2I�S � DSe`2D     ��� �����*� ����Z�Y��Ƃ������&�����b��n��c����ߓ�� �߀0(����/��������6���  @ ���?�����&�(?ԕ�  ��������  1���É�����	���j��ɀ 0 ���"��b�훤�J����?��ܟj �	��c�k      �\�ƴ ���K���/_�'�P�o� ������� ������2c�����C�-H��N%�PE	�S� @��2��s����r�v�6�ɀ ��� ����ݳTT RQ��D��c��f���J>

�� �ٔլ�ھJ۠/������)۠N���٬c� �   	ct�۫��3]Sa �	+ � V��	�?����']Pl���������iߴ������i ��c�g��w��7� �����!>@/�
�� ?��
�J�
� /�	�
	&� ���É� ��� �������"��� ���c�����/﹛ ��&��������Ɉ ��c�/ل��/���k��'� �!.�/����F8��;��oy;]���~ۍē�D�1L��                                                                                                                                                                                                