��� @d @ �� 			     }:> 
    ?<"~ .���������                                                                                                                                                                                                                                                                                                                   ���.!nEfFb!�⨎������㠕��.&X��і��&ѝ(� �����㠲���&��2@�␰���0��'��J�/�è��ϝø� �Ñ����� �   ��6��&��C/�d�0&0�1�j/?01r/�/ N0�J���i��bi ��Xp@��u@ee�@ BP���@�8� H$����O> ����!H�.!.I.d�&�/&��0cH��10b��ϰ/������6�?/(/����l/6�6C0�l�1&��� 0D0�	&1�)87f�.�	�y	6r	�{ 8q.�.n7!.--&�a..�.-�/�E�F�i��+ ��o0�?�d�0G&GE6GGCF�l�Ւ�ض� /��@� � N� ;؅@� �	
�⎶HD.!.J b�!. !b�!.!"b�!."#b�!.#�i bD �..&...bgw �J��ï�c��/(/����l/6�6263646060D.0."	�l2	'3	'4	'�"�DD�..&.&!D.!."..b#bDD�..&.&�����c��/(/����h/60656� ����!�z��"���H�!5�)1&1D>12	6b!1�1@...&��.�"���..�	��	�6	'.	&5!.����<	1t�0���{.&&)(/�@�..&��.�"���.&.&�&��(��/c��b�/b�l//6�<�|/�J�F�E�i��+EFf����׳  ku�C)t&(?���G�s �<m);�&N�C��dr"qH$�ؤ"�/���b	�l/6(?�.0c(��1�18&7�lZ/ਟ�0�)�1�08&��)�.�	�y	0r	1r	t"�J#�/���b	�l(?�.1c(��01b87f�0�����.�	�y	6r	1r	t#D��� ?����  ���B��b?�l�<��K �|ly���a�S ��O�@t�sH�A�
�%A.8n$7&�.�-bbKbF���'%q.9n$!.:&b�&r��r@,b��� ?�a.�.�!>+�/��"L�i/�b/� ���/� J���/b�/�0���0�0;0d0@>�,<n;"F�/�L9�:�<//L)9�J:�J� ����ߋL�ߛ��d�����3���  $���  �V�4{ ��\��CD�����/������%q.9n$!.:�g��?� .?&b��y�9��:���F��&IK"���H�"������õ&KJ"0Kbb	�l	?0t�Ш� �K�J��b��&�/K�|� � -F���+��� ��&�	&�/&	7/�J�־�H>������?�/"� ���(�?0B���@��p΀��� V�\ 1h�4��?�(���i� P �
�����F�i��"�����r��y*(/���� �   ��� CBAf�D&���8�BB&7�AH.ABbB�C.CDd�B�7Cb8�k @˟��Մ��&�@&��,Ё|��K   ���   �ѫ ADA��D&AP.�@/�.D�J�66b�r����$� ���� �������χ� ��� ��i�����,��|��<�������<���'�!����7�����s�Θ��'H.����~� ~��r�b		c�t�'�-�k�����J~�)�Ê��&��B��ry�/4@�~����� �=kR��b��b�@n�u�N�*u��� �M�/|���c�V��y����J���P��5���U �`����+Nd !������g�'�'�'�!.D�/b�a//������00!.H/�/0b/r����u��䎶��r�s �����  �����r��r��r�b	c	�t����������� ���>�����0��&����������J����P���/�󩀀�׈/� ��������]t 8� �,��&�Ά!���� �//c(��J
�
��/�8/�J��(��(���� 1��   �� ��(� �!��&�Υ ���<��|��D��J���  /t�b��bj�gd�2b�� �"(����/�ؾ�|�2�J&b�bbb�j!.�/�a�d����w����w� pp (��n')�H��T�?  
 �o ���(� ����(��ϖ��E�,��c�����8��(��(��� ���F�(?�����J   !��&�Χ ��������.���.� ��������(ĲJ� � � �  DD�%b#%D ��#&|E��#�b�#&##6#e��|��*C^�/��|i�a�c�� �khPoH���4#�0p
 F E? �� �� �� �� �� �� �� �� Ԡ �� ��  � �� �� �� �� �� �� �� �� � �� �  �� � �� �� �� �� �  �� � �� �� �� �� �� � �� �� �� ��  � �� �� �� �� �� �� � �� �� ��  � �� �� �� �� �� � �� Ӻ  ��ז                                                                                                                                                                                                �����2����&�	&�ǁ����	(?��������   �	��.�ǁ��	�Z�����	�A �E �5��9��= � �  Pց@��@ց0��@F�P� 4֌@� 1� @��0H
� ��������ׁl� >��b�8p� ?��"�����'��J�����+_ ���߄������ ���)����d�߉����w��s������   ���Ғ������?�Ӣ������l��6����b�|��'�J�������2@�␸���0��'ޮJ�.T���>�����0��&������DƁ���,�Ԟ                 � � �����
G�JO� �
��� � 0� ���@80�I� �������� ���&��6�J>

����� ��(����������(��(� �&!̟���'�0C�LN��P5S�@S���8NXT "���Se`2�3�NBՆACE"�8�@1��DM��C F�@)�2��G��@)G;�DH+   ������� �� �       ����� �E� 
��P��
�  ?"                                                                                                                                                                                                