����   @ @a.3      > +
0&0!+0"+66#62> .?      : 61</%++4'3&"'2/    _2 :  !!!
0 ?<`   : ?>( .   00=; 
" <*3'>'=<> *-';':                                                                                                                                                                                                �
 @ٔ�MA   �!��3T8     Uo#�X33�1  #��!�!������۪��"��$��D      5����  ݏ� �����                                  �    ���  `             i              g2�� ��`���f��?��X�X="�o �*�*'�%*I'6�?G&\Hf*'�OHB7)5)_H"Ii���\�NIHtG�J*'�VI���\!.(��\[i\.&.E&MhbNNc���NMD��M0 D@�M1 �6�Pi�B�C4bDi�����B3"B�oCDD�E��.�EMfhN&N�?�N�M�JM�0D@Mb1�6P&��BCf4D&���} �.�����B�3B&�C�D�JE�K8 ���q�K*'�*I']������ ���&*�*��2��o�'i*�'���()�D>���'i�O2(���'i�P2��(���b�b��n�b@��D����$��F'�(9�O*���D����D�J �P     �#��3��?�naih �    � �� ��  �Oi9J&K:bLKb<B+PrC@",,s�X�")P&)�-�#+�$!�� �8�/�K�L�OKKdJ�J��K����*'��9���� � ����R�R�+ UUT&U�-���� �SSb����Κ Q��y���Q�-���� �����ޚ ���� ������ �-&�Y&Yt�� �������2�ޡ��x 9JKf:L&��^-b#C�@X""P�&��K< B$)!�� 8����R�!���^Qb2P!,㨮�,V6Q2 O�j+!>S�/�U�SO&+V6�^����K0"KLd��������j��6�O� ���*'� I�Ϊ� ��/���2 Gb���_�GG&�G��\�WG� G�_H"I\d�I�HGD�\�!\�W��n�2��" FF.
2�7)F2 7)� �����������  �>b��b27��d�Ѣ�� ���4��c�(�@��

�
��0(���@/��"��������@�� &!��"��ʠ��?��� p����&�!���6AAb��u������"�A!.��/�״A!.��/��K� �U	�����w �%@�X")P&)�O��%�!�� ג(��נ/�%�6Q""!�� �8�/���%�����*y'�������.�(]�.Ng� �������ː��b��b��c��c��ɀtͿJ� ���   �P�����ź�  �8 �����6Z�J�Z&��J���d� ����@  ��=�&������@��$� 0�26 �������6�=�b����P�   �&�	&?�&	7��J�_�h  �NĀX�̀ԀN���D���D@��TR��	A�HT` R���ET`!�T@SX��C ��	�T `�TS��� 0`VX�A3 �TE8LNb�GI � 0`VXCLB�$XM`	���N�/`VX� M�`�	�3R�N������ #	�҃A5RS��P5 ���� #	�҃A5R��AM  ��L USA	�S�H��5�`F��E�d�8҃� ��T@S��  R`O`eՅD���T@M�`	�J`G�I� ��;�/A��!@�������}R��_�����Ȁ�                                                                                                                                                                                                 �����������������I�+���)�����������K ����� .��d��J��d� �    �A �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ޓ�(��@����)��J   ���� ���&��'߮�����w��@ �?p����p��w� q x ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    ��}oto�nm�{|� ���f��f� g��r��������i�����g��π�ܠ/����&��I������   � >��y������������c�� �k�:�ew�w@�����wST� R���������6��H��h� �   ��)��9��� ��?�>��� �������)����������TN"�  �	���/���g��)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP�����w ��:fC hRT�S����wހ F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�旓�� � 5R���D�� � �Cv�g: hST�R���� � �� ��� �����A�����рh�����������=��E���)�H���)�K���)�N���)��������������������y������A ��LD!  ��N C�� �Q�> ����������� �tq� .&�jK)����&�J��' ��&~a.i�6��ik9i�2� �O�wC�g 2 q                                                                                                                                                                                                