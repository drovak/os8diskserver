����  �,%  	#<
: ( *"$  *  ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                     �+&@ٔ�MA�� ���L �Z�I�~�� ��~� ��~�����~� ��-%J�~�%� �F��.�{&z�'x�'3���3�������� �%�������������������� 2�K��� ��\ ��I?"�� ԅ����6�W͵�[% D CP�(��� � � �@ ����c��b

�
�菐(� � � (��@/������ ����*� /������&!̥���?����������  㸹k � �������0�c����0��bJ��
.���d�ジ�r���"�d�䂸�r��d� �    0����� u (��|u |)�ظ� �� �(?��� ��8 �����r��r��y��������������ْ������� ������� ���������􉝁�� �� ��� �� ������~�}��� ���Z��Z��Z�������~���� �����������~�}��������咭�ꛀ���� ����" ���؝���۽����������~��݅ ������������ߎ��� ����� � �������-���(�������� �������w�������������� ��������}��ڎ �� ����٨����J�ъ���ǀ������5� ���J�
>

�堮��c��@��b���� /��@� �P? ?`��� �� �k�"��������煒݇����?��� �������� ����������(?��������}����Z��������}��ږ��������&���ܒ������������& ������݄���� �����~��9�@�ؖ���s!��(������ ����Ub!�l� "@��ْ� � d ek������"������'��~��s �n��~� r��݈������� @���s!���(?������(�������'��������݀������w��=���� ^����!>�(?����(�������'��� ���� 9�����4(���/�פ�ף  kq�s)p&(?���A�o � �<��� @,�������� "�� ������'��~��=�������s!������2��Z��������w����'��'��҅�ݧ����U�����'��}����^�?��'��' ���=��ڈ���!>� ?����>�����Z؀���7�ʚ뮺r��  ���?�+ ���Kr�������w��������� ��@� ����y����"��J������&� ������~��&�����������9���ߟ����Z���� >��&�����������9��'�����������������������J� � �c�t�ʫM������ݢ�!|�ԫ�����d��6� �   �ۢ�݂��d͊���  ��� ���d��  P !Xπ����_�"�. �����'��'��'��'� &��w����������r��r��r��y����넟������� �	�����������) �	����8������)�����U������)�	���������&����ф�� ���㕉��� �B1��������z��D �a��bD�5����D�� ��c�W ���"� ����� ��������'�&�&�������󙥥����������������څ� ����w��U�� ���� ��_������P 0 ������@� P�� ` .����^&����T.!�	�� @^+���E�4^&���S��&����� �����U��UU �U `����ـ�D w��X��!�� ���Z�����F
��!�� ���Z������D>���s��7��7��3!�� �� ^��Z�������s��Z��y��w��s!��@������Z��~��2��s�@���������!�&�d�&���%2%+d�%�] ?��� `!��k \������� ֈ�������U��U���b��b��b��b��t��D�����y��&��&� .� ?����J��J� �      ����_����}�����}�é� �n��~� r��� ������ �-��������ZǄ������Z� ��������c��������������J��#�����Z!�.�Q�Dԉ����������ރ��� ���� "���&�&��f&!̋&��ď椏�!�ʀ����f@�����J��b!����f�����&�����&���J�����&�@���"�o�N��b �����!��������b��n��"��b�@���o��̀��+����&��  �          �	��f��f��f��f� u �U���k������ ���)��)��������)��)��������)��)��������)��)�������)��)	����
���)��)�������)��)�������)��)�����0= �� ���i#�� �  U= � �@
	  �  � @ 7+ � ����)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��)��) �� ������������������������������������������������ě�Ĉ�� �.@X�
��R���@ �� @Q7D�+ � ����'��'��=��ْ�ڀ ���r��r��s��������������'�	&�
&��&�	��
s��s!������J� � ���'�(�񒍚�� ����� ����  �������ŋF��ƴ����� �P (����DD�����DQ��DR� @����C��O � ��D����݊���� ����߀�� ����) �	��)8����)8����)U�Y��)w����)��	��)<�������)�	��)��������=����@����������=�����H����������s������@�ʀ��Ѻ���=������H�؀�� �                   :	��w @���}��w�<��S �ǡ8����   �����n��b��b��ـ�⁇J�������'��'��=��ڒ ������'��7� �@����Z��� H�󥫝�� �@����Z� ������s�Z��~����!����5�������ۘ�����&!���c��` 0 N�`	ES`����C�$C���K � �
�4�W����P҈����@��������)��������)��y��������������������}�����=��������ـ�㍀���)�����������򖚶��������@����������+�������0�����W��������"��c��c�ݺ����}��������������������Кz�����wŋ}8D�5z�� ���&�"
�: � �D�̀���D>����s�������r	�n�	���Z�������Ũ����ň������b��������s��������������������>�����8�ś��8�śF���ٺ �g����� �-  �����٫ PC  �^F����Q�D7�+�� ���݀�� ۀ����'�	&�	���Z�����x��7��B��r	�n�	7�	7��Z� ���r��j��������&�v������&!̱�� ���w��'��&����7��4�����#�����Z�������&�������J����^F��   �^F��ӀL�^F��:��@����������� �������ވ������������y�_���'��'��'��=��"��r�����r��s��ّ����� �������Ԗ�Ֆ�������r���ԅ-���r��r���ԃ-�뀞�!.֨/���J��ֲ��r��y� � �   �����"����c�00� ���  �͕���Ԫ��� }6�����������5D�����.�(?���(���������'�����2��z�����"��z�����7 ����r��s��Ӆ�ݧ ������'��=��=��� ������	�߄�����~��r��s��٠����'�=��!>� ?���s��!�� ���.���xTӎ.��rÎ:	ـ�-6�����>���������� X� ����ɀ�����c0�0 �������� �00� ��������������������c�0\ �� 00 ����������c�0L ������� �"���'��~�&�&�&��� ��ώ� ����� ��!��"���&<����Z��&��B� [��   ���8\  ��ڱ���� �@�Q	��� �	��c�00� �	���ɔ��� ԁ 0�0� 0\0 ������� �()��c�00� �	�7�8�ɕ;�<�� ā 0�0� 00 ���������ST����NO��c�� 00�N��00 ���������de��c��� 800� �	�ճ��@1�N�� 5�N ��`1������Q	���_�����0��2��y����@~�>�~��s

�
���>�>��s���D�����c�00� 󉆾ܾ�Ʌ����ɖ����ɕ�������0�`00� 00� 00 �����Μ����c�00� �	�����ɑ����� �� 0�0�`00 ��Λ �D��� ����:�Ђб�w�Q� �	����c��T@��  ����!�� ���ҕT@!����D@ ��


���s@���s���>��y�9�9�م<�=�� ��`��0,`�00� ���8��ic�0 �����ӆ� �� 1�80< ���8��i � 0<�� �@�������p�q��� 0�� �������������p�Q�                                          ���f��f�(/�@��/�פ���(���H/�ؤ���(���H/�٤���(����$ �����֜d�F.���"��t�F.���"֜{       � �� �� ˠ �� �� �� �� ԍ ��   y ����� ��0��
�d��< �*�*��� � � �=��}�Wy���C�iȥ�h�O�h�`i楇���K    �fb�2ǲ3'4'�� ���n�[b�!i�� �3�<*)���D�懺J�� �����b��b��c��cߤ��t��J������c��m�dX̃���NĀҀԀN�̀�D��C��T@ GS�TR���@MN0 ���R��C 	�H��HGS�TR��AX�K@��� 0�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C C G�S%�RA��D�NS��S!�D�H�4T@�����7��� ����    {�������∇r��{��+�����DD D"'D+5D��D��D��D�EUHJUPRU��U��U��U��U��UԆW��w��w��w��w�.xJL����������"�, ���wLN��`�b���������������ę�ʙ����H�49 ;B DF ါ         ((�  pp�pp�pp�p(�$  >                                                                                                                                                                                                