����  �
*8 
>? *	$'"/<*   : *%00**'8 	!>? *$'#"/<*  "5$',./  $=#?<559 <+	+: 	 $;; + .50>?6??      >><8!>9888!'$?                                                                                                                                                                                                 
  � `:" � ���/       � �'   2gFOw_kw� xBH����ڎ��( �"��"��"�c"e� ��" 
3Q1K^ #IO""	�   � �                                  ������ �����0� U�   � 0���U�@ �H�@?�X�/ ������~`/���}"KKc�<i �K�<K�L�==�|�D{bz�{ ���O�h>�M�>�!N�M�O.���'p����>���O���>����� ��O�NOdOK&OOBMKcO�k 	(�!�� �>���N����f�h���n �bD�.Hs�b �J��"�*n &��,�m� ��K6��CK�t� ���P�kFQQd�P���� V&��V�/��!��"VƖ ��E� ���⾠/�����bD��濾#��r���Fʧ+IcAc��aG����>�.   |�!�� ���c!��ѠO�Ѥ�ݲ� � ���6��C��d��6ހN��7��D��J� �   u��#��r���"�a� ���6�'I�����
    ���6d�
>

������� �y� /���(�����K��b!(�����x�&��(w�&� �vH/ut";��    �	��� ���sΛ ��C!��"�VCk'A����., �C
�C��n�bQF�u�7� �P(/i �Oy��m�L#� ٔC ���6��C��dr�!J
�
��rB �ᔀ� ��.q�q p�'� �    ��6��K *	9*N�<�3�'y6�4�(?���' �>o���>n���>u������K> 0���R�d� ����S�d� �>m����>l���:� B�� �9 ����Y�*e��*9Y�) ���;����A&(?�6���� 	�ʀ
� �̉�� =	��/���ʗ�J� � �@��=��Q�>��8�SD��� �� �      ����⩩b����k � �����⫫b����k � �6-�H-iI-iJ5i�ɫ =	� .=���7� H� ��7 �I(��؂��7� J� ����K��J� � ��P� !��&��<���k ��<i013�����k ���&� .��b���� .���!kఱb� ���⳵b �浨/��� ��!.k���+         
 � � �  �  � 
 ��Ca QN%�PE.P      ?	 	 
 ��D @ 
�DA @�� 
  Ɂ��3��@�L�C.� �  � ��� H � 
 ل�MA�Ŵ 	UE8LY΃�N@ NR��
 ��A�EG�S2��3���	�NB�V&r�B��>�bWr�c�t�ʫM�� ��ݢ�!|�ԫ�����d��6� � @ �ۢ�݂��d͊���  �������J� ��w)  J
�
��(��H���=�=IE���� ?8�A�B�	��R�J)�  ��A���B��4?�	̣	��R���) � �
	̯	����E?�
	��)�  ��	����R�J���B�b^l�]�]�J^�J�\&��	������J)�  ���	��	��� �\�J� �                      �� � ��� ��ϐ���) � �
B���                                                                                                                                                            ?�	̅
�	��) � �
	̏
�	�ʑR����?�	̝�	��) � �
B�	�ʧR���                                                                                                                           �?�	̅��
�ƞ�/�R���*���*9��S) ���:�
� �  �=Y�"�
� ���)`� �
�?�=	��	�� �)ɠ  �=��	��� ���R���	��?�8��A�	��B�B�	��)`� �
���	��R�J)��  �A����B�	��� A	,B�� �A�B��=�=iE���� ?�̗)�  ����ʔR���3?�A���B���R�J)�  ������ʰ�M?i��̹���) � �
������ƪR�J���b�b^l�]�]�J^�J�\&��������J)�  �����	��� �\�J�\&\�J\�J�@� ����� ��ϐ���) � �
B����?������R�J��?i��j,��R�J� ?y��i,��R�JӰ����̬����Π���ō�������Ҡ����É��������Š�����͠���̠������Ġ���ȍ�������נ�Ҡ��Ġ����������Š��Ġ�=�|"
�� �)�`  ���?�=�.�~��� �)ɠ  �=�-���� Ϊ��R�J�=E�04?��3S�72�-1��S��s��R����0/�6h�E7i.s��6�=E� 72-y ���7�2-y1 ��0�/<���"�h�E+i.s��<���"�=�E ,2�- ����,2�-1� �����=E�0=D? 6[�=��=Δ=ɑ��x��ZZBg�/�����W�/CZ�f�/C�WCK 8	�Φ ��
�YZbeZ&Z�/�W������Y�/C=���?����72�Y1)C�RCK=ɑ�C{�Y�H=i��C��YI&=ɑ�C{�Y�J5i�?��=���C����Š����°������ҍ�������ٍ���΍�=��=��=ɑ8=�= .dz'E�h ��!�k�/�������*�*��*<���:*=���:) ���:�  A���B�	ϸ'�>��
�Ƽ�+     �k�����=E�=�k.	s��.s��ţ���٠�Ơ��̠��Š����Ӡ���Š������͠�ӭ��������Ҡ���٩��������Ҡ��ˀS�D��c�b�&��	��R�JS N�R&����'�Z�8�� �S�j̟R��S� a�R�o���'c���� ��S�'l�� �=٘���õc��F��6�@n��"����F����`";����D����,���� �   ���|!�o_F�!��? �	��R��B�� �                        