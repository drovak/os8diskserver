����   � �?   ?  	!    ,  	  !  	    !                                                                                                                                                                                                                                                                                                y�2 R               ��� � î "3?"��!!�  �                                                                  b� +$                              �70 �                  �90��ǩ2 � �����������������Ië���)�����������K ����� .��d��J��d� �    ��@ �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ޓ�(��@����)��J   ���� ���&��'� �       �@ �?p?�/=� !�  !�� ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}to�nm�{|� i_@IQe���r��������i�����g���ˀ��������d������� � � ���������y�����y��� �����Q�!@�?>="��"��"��������6��H��h� �   ��)��9��� ��?�>��� ������������������TN"�  �	���/�����)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP���3>"  M�À��"�"=?"�  F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�f���� � 5R�� @         �� �����"� �� � �� ��� �����A������l���Ήl����������������)��"�����"�����"�����"��������������������'����� �ρl�'��6ς,� �   �� �LD  �� �C� Q�� 茀������            �   K	��� �   ��L 1�
  fL3     8@ �    nSl߀5�FS U��50D̀4�*6 �E�a%�bhlUp(3    � �� �@ ���?���?� ������ �                                       ���� p���R_wJ p                  �bf   Y n����n�� �~C��o�&�&�&�&�&?I&��7�j�gI�Jo�k/-��-i�i8�
� c��I�GJ&0IblK&-Ֆ�-��7bI%)8%)$��Ī0�NKItJ�J0�/�-��$i˚���-�$����8�
D�ppbc�/���-y$y�������w�v�d� � zKq�5R��8Tqi�r����-�$������
���t�n�-y$y������D�s�8��s�stb���p�/54"`s☕����-���'$��˪��'EI&�i�/i��It��o-i$y˚��� ��/��K 	���̺���@� SS�-�~�RH.�����~� ��~�rR��1��|}w{�p�����?�p����c�/� �(�^�^c"ș�c .^�c� �t ^^&^ ��DJ&J!.L^b�54"I�c� �sI ggb I�JI$�W� V�^ ���f`.V�/�W�!V��/�f�ViF�_i�oaiIIb	@~Ia"�aOdׁ�u�/���x  ����K                  �' |'}zwMMB��MJ.1RM2 D^�^�c� �q1 ^^&��? r�T�c���^.���eT"���T .T!i ���u�"_������鰢yufF_&F`&m!i ��m��Ԛ`�J�Q�5(�n�m�I���uom_d�u�mnf�u����y�JD�ȳ�_�/�u������S�#�� 	���h��@�h�i���X� (e��1�{ ��b�Sb3x�2b��Jk�&n�/������U6 !Y⠩��m�(��H�/��C A�A���7�AB��_�yF������?�/�/������-�݀c�P&P�6�-���-Ö/��P�d��6�zB��bEb��b@��D����O/����D��n-�.9��JPF2�{��{���D�,�D���d�D� �O     ��/��f��f ���c�k ��%)�%)%����  ��F�&�4 7%)�.�樜J�� �/����F���?(�@��

�
%�B0(���@/<)��J��� �%ƛ�� ���6�B����̴���r�r��r��r���    	��� �;Q&�I�6JUxb���|S&녵���   n���b!.a�/��&Sr�D"JJb ���b�"X���J�&T�&�� Z�b6Y\�	�]�	[&]!.\�/�b��n��`�&I���J� NJ�&O�J&�?m&e�~�& � �
   �����"�n��"��&����"��b� �����F.��b
����b� ���&��&� ���&��&񜲸 � ��Ѹ�� �����& �����,��u��<� ��&,!��"��  ��b��b�!N��/����!N��/�����  4 l�&��?��K 	�� ���'�����'4 Ib����0IblI&�I��I� J�IIblK&�K�I0DJ�J
.4D �c�d��K� � 	����M4 �����P(�i�0>=" �xnfV*)WX&TI&T@ J^b�)9S="|Ib6J+��bv��x�/����O�!X�(��!}�}!.OO&S����	}t���b@.	?}�b��O¨�������K���I NLX"X�m; /�X����x|b�I�6J�w�Hv�� ��S�/��_b& ���������J � �~����xwbHv� � kSaf $	�c47a�␖��0H
�7 .�/��4���K F��f8����O���ꘘK M4��j"��ng�#�� �� y�@~�"��e�d2�����r ���2"��J��n�_�/y-?�M4 7%)�-�By������� ���~Q�Q�+ �� UU�-�~�a�~-�-�<-)'�� �a��3 ���
?N�K�EbN�ni
&��+ ����)��&�!��"�ΐ ���-?�M4 ��b7%)�-�%�y�l"��g�Fb��b�������J/-�?�~--�~ �!W�O�nV	&o�/�E�N�ni
&^ C�&��+� �9��I&�J&IK6K:0�K7IJD��������T��D�lA�qoiUbeQ��b  	�/�-��G�&��f�2"��bk�&�)�/���7%)���.9��D�����J� �       3 �?b��d�᤯��)֞,(��'�@��>��,��")(��'�;�/���&�@/�/-�|i� ���K��K~ �������    -	�Yb.��-��Z.)�-�[b.��-��\.)�-�]b.⛅�@	�0T`R��	A��C��0@����X����A������倗�S����D���စ�DU��ET`!�T@S P��@	�0T`�T@S P	�T�@��C ���� #L�A� 	5 XR�� @S���#��4υ��@` X�D1׋M��h6-���C��ă ��$ƃ �PP 0�L? CP�  X`���� @���#�5���_R`O`eՅD��S� �C1!Q ��MA� Q� [�8S�"����C 	� HS���@P3@X                                                                              )}�                                                                                                                                                                                                