����  � �� %8.6 6 7 7 8 8 9 9 )��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                             
 @`�MA�� ���L �                                                                                      0@ � ��  #�����������
�6��U��$eD j2
rl"C�"3'"	)��A� m� �tR���"��"��#P�t���k!��/�.�������u)�u)��(����u.�H .)Pn)�)�) !D�)"�jt͜ �o��xik!��/�.������.!.�(/������u)��� (/�Ы��.J 
�
�wk������.H wik����/�.��Iwi� ��� �� �� P �(?�r�� ,
k!��/�.�!�⨙�.!.�/����&�u)�u)�ߢ&�u)�u)Ru)k��/�.��Nwik��/�.�FZ���..�Swik��/�.�FZ���..L�&k!�R /��r tt�ݵ�� � �� �� �P �#�"��i�� 323F]3��3 �D         h����!"f!6!!Cb�J�#o��)$ti�#�RK"uw�"q)w$�q��%�i$�O��Z�#�/�I�&!.L�/��L�
����O"b!S⠕�S �o
���K"b!O⠕�N �oI���F !F⠕�F �oM���I ���H �oK��� I�bI! /�!�""B! ⠉����� �	7
�J� ��	�
t��� �.�Wb
�o%��&	6� �n`�a��l���&沧{� @����&� ����BH��׳�   ���H�� γ���K��b(�ר� �� ���F��b@
�
�S&�/T"�k ��&!��.�.�+�<"�i;)�f��H/ �H bI� bFS&��bNS bL� � � /�n�j<�(��l����Knj�E(/�l���������&� ����I�� �ʠ�̭ˠ��K� �-� ���,� ���� ��,��-�� ����ӽ�� ������� �yA�N!�8D�EA; x	�2�r�� 71� �foa�ge�`l���� �O&oinj�< /�g�ei�l��m��� ��Q�fon�j<� ��ge�il��m���� �Tboigj�e`�l��j��89fdl���� �O&T&on�jg��<� ��ec�di�lΚm͚� ��Q�Tboing�j��< /�e�cd�il��m��ݫ��&�@���E��� 0�H> �O&T&on�gj��<� ��ei�l��j��E(/ci�l��j��E(/di�l��m��� ��Q�Tboing�j��< /�e�il��j��E�(c�il��j��E�(d�il��m���� ���'��'����Ձl�&��t��� �� �xy�^T�`�	B0LT"`�m�Rxx���
��(��H��� ��/�O�Q�Tboign�j8�>9b?iil���&�nj��<⠩�>'&?(&e��'>&(?&il����&(/�j�<(/�l��n�jE�(c�il��n�jE����:!.8�/�;�!9���:'&;(&�/�8�:9b;:d;�d��':&(;&il��j��:�!8� ��;!.9�/�l��m�����R�����@L@@F��D o	T&Q&���e��& /f��8�&9�&8b!H� g��&�nj�E /�8��:&9�";iil��nj�E /�:�';b(b���8:&9;&:O;dI�'�:(b;iil��m��n�j��8!.:�/�9�!;�&�lȚ�&� ��m��� �   i��� n	jߒ(��t��t������(��t�t�����l��䫵�DP鄣�S&��`i���J�f��ai%oge��/�c�d̝I���� ����8�/�9����%�/����)T bSK �]�(^�!�bM���F���bb]�/��!�=&F.�&8>&9?&�_���Xr�k��R  �ߴ��
{�/�{��&,���   ���7-� ��-�խ��݅խ�-=�-[�-�&��-Y"����Ι ��}Y�����I�/��7���&0XBb ��I"�f��Q����I"�f����_P� *�G*"���U)&)�J*�J�˺�/��I�/g˛zb�I"�/�����t��sw�=!.q��T��� ��X&�IРb����@ � "b���"7�    ��&��Ȧ�����-�խ��ݏխ�-=�-[�-�&��-�Ο �!}i|,�ȩ�X&�{����t��s�t"�,I ����-����~�|��,d J@y@�� 89��(��==&=^"���].=�/��Q(�ܻlR=&f�*�8���ת�x�f&x�8xkBfxc�i�i�J� �U�� �� ���� �8�/�9����@&Z+&Ҍڀ����Ԓڀ���-@�-[�-�&�-�Σ ��}i|,�H��I��� ��h��8!.: /�9�!;� ���K� ��h��8!.: /�9�!;� ��� �_P� *�*G"���U)&)�J*�J�{��Q��,�J���t�@��t0�sw�@!.q���v�������� ��� 7F+"���,J.��M��B�A�D�Nh��O(���Z+&,I  ��8!.:�/�9�!;�(������+d�C����ʨ��W� �@�&8O9B(��@@&@^"���].@�/��@�k ��խ����-��-~ʛ@ �� ��@&�8�88b���9� ��8�k�9&�<����� ���b ����+ �
��?�. ��                                                                                                                                                                                                �,   ��@�.��                                 ��"   LG�2                                  ��"� P�D ���2 @����ͻ                                                                        8O9tI����<�l� �
.
��t �/q)Y&/�	&

d	6(/�x�t�
v)w�q
��J7(/�t�7�q��ht�Otɑ����� H��tX�Dq)t��Cq)t��Bq)t��Aq)�E� �                                                                   J)b�vw�v)w�
�v�F��)���(8r)9

�F������"�  � `�ti ��������������л�� �.�Wb	g	�J� ��p�wΝpw��p�wɝpw��p�w8�r9�� ��8�:9b;>b8?b98b���9�/�`��ҽ�խ:!.8�-�-�����-~՛@<�� �!���� .! ���6��6��&��&��C��F��4�@n��"�n��"����F��&�����"u����J������             �����Ϝ��������7��ʸ��Ш������U�ҭ�խ��-�-�����-~���@��խ�����-~ڛ �/@<� �瀮�-����̭���������խ�@�J���s� �����"��k��_�'-�Ȑ�?*�g��1�� �C���A���*U�R��� 
�
'	�J��������*@��(����f�F���h'	�J����� ���_io����������	tŀ�����(�b����������}~�� @���
���
Yb
c	t���J�?�� � �!�A �ǁ0MâY��8�
&
'
P.@@�	�ǫ ��	&[&������@��
&Y&
>��b	t���J��� b�	t��'�y������{���}��Ѐ���"�����&�D.���b��7�.��4��b��c��c���G�O�>� P?����@�(Rxp@   ���6 ����� ���b�Ȃ

�
���
.��ț(� �H�u�� �Ru)Ru)Ru)� ���f��&ô&��@���/�O�����"u��ɴdʳJ�Ĳ�����    ? �� �� ��� ��&�6�
.

�����֊   �(в@���/Ru)� �&��!��"�� ��u)�u)����� x	yҕT`!�T@SX��C ��ɀ �xy�N �8P@���� y	 2�0 �� �y �5v� � y	 8�0 �� �y�� D � y	Ԅ  @� �y��`3 � y	 1��IÀ�; y	 2�0 �A 6� �y �10� I�5X� � y	 1�0 �A 6XN  �?����� �k�]O"�62 x	yҕT`!R��@O� �y��υ� AT � �xy��DNN �P �� y	R���T%� =	ES��K x	y��DU�RA��D����� x	y��DT` R��O���� �xy��D@S���K x	y��D��C� @�`� �� 5N���@1�N�� 5�N ��`1��	�8 x	y����4υ��@} � �xy�����4 � x	y�X��4TS@�� x	yϐD8N�P��4TS��� ՁC�N� x)� �xy��C���E� @� �xy��C�S x	y� T T�A��4��E��4��; y	��2 � x	y�� H� �xy��TR`P 0����߀[�À� x	y��DM T� �xy�� E�D�O1C��1N�� x��������  �@`�� Q�$ �D��U �#� 0�D�C��3�O��8DVC@��5DC�TɅR��C��R�� 8�(�� ��TO�#� DT � � 0�� �   �P����� D                                                                                                                                                                                                