����     A('  7+(7*,+ T :6>(*?7>(*:7$> .: 
./
 ./1!  8>(*+?7<: 7:8 
0>(*);7<: 7>? .:
../
-./
?  
7"9
8"9.1
  0&0!*;: .9  0+ 0>0&0!+=<(/<;<(/:9<(?8                                                                                                                                                                                                �@ٔ�MA�� ���     �� �� ��������?D0   �&���(��#d�� ��8@��7��@� ���Ѝ� �   W��?���� ?V������������� 2�K���Z֩A�?�����s�
��� �v���? ���?���R��`����ȶ�@�JA�J���!B���&�(?�B�����Ĵ�6��C��d�!>C�c��t�CD�����6��/@�����"��j      ��2�����2�����&��C(���������C�F�۵d��0��&��C����b� ��!��� 
.

������ u (��|u |�/?��� �yW� �S�_�Ql�l���	 �Q����  	��A���� �Oj��jd v�O"�p
�
��� H  �y |���D�PQU��A	 �o ��D" ��P ��T                           �$b	���F�H� ���@� �����������'��'��-������ڭ���������  �  ���������(��������t�ګ �B�������������K����?� a� � ��݀�����ꮻD� ���J�
>

�堮��c��@��b���� /��@�v��?�?`��؇��� � ������� N�������� �H/��O�������j8�   ���ƌ�+	������!����̯�&�����"��hˍ���&��&�톖����ގ���"��* ���O� ��F.���+��   	���F�H��	�������j �
'�	a� �����᠎��&��(���������္���� ������	��F
�������h�� ̅ � ���� ��)��)��)������y�zzr{�}��݂�چ����"���Äڴ�툉���r�������>���D����߯o�1&"01�1����++���,�(�1�-1& 0&�+(d' ����+��� �9ŋ�N��ߎ��ڨߑ���ߓ����+��B���a������-��� �⨩�����������⯭����P� �(��(����  &!̻��� �����&!����(���(/���(���� � ���-�����'Ӌ���	  ��.@V ~
 � ����� ���?r ��_���8 ��)��)�����������F����������y�����������(��
�����ڎ�҇����� �������                                                                                              � �?�1�� 9�P