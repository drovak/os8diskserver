����   H � -       --      	         #            .  .   ?   ""   	 	        		 =  	      0        	                                                                                                                                                                                                      �                                                                                                                                                            ���' �� t CS�����?�����p��n��c �l[Ϛ!�������������, �O N��É�Ϩ�� �� O N���   �� �� ύ �� �  ����"&�#&��5$���� ΃�                                                                        >�&3�  �'⠬�&�/�"�!#⨬�%�/�#��#d#�"����#&�����/�'��ʢ��/���&'f�ʢ&��$�k����*�!(⨻�(�6�~ ((t�'����'�j�$�"��&&4(&�ʘj    �  �  �  �  �  �   �  �  �  �  �  �  �  �  �  �,   �  �  �  �P(0�� ![��@h~�(��}&�"(��� /�%���� ��%�k�(/���(��� /���&�b#�b"�j� /��)�b*�b&+f*(&��(���(/���+�B�n*'*�B�*�!)⨧�$�/���)!.*�/�*�|�/�{�*�n**&*~0�(/���*}0���*(&�*ܤP*0��u��B����M ��� L !�� �+�/���������n,�/���������� ���� �))4~}�b)�/���)b��������6,�N�+�n+H/+�,�j ���6����l�(/���z���&���
>

������ �y(�x�H����&�ۛ��� �       �  �  �  �  ��� @ 
�&�B�� ��"7""B��/���#�/���""b #⨏�$�/�$�&�� ������d��6��&��&��&�@n��#�n��#H����d����!>��&�w"�ϓ� O�͔��D��C������          �  �  � �   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �>�"��3��i@i� ���ƭ�/���e�������f��#H����J!��!�� /��b���w�"�����㠎��w"���i��� �    ���   �����<����<�������>����< ���@�!�i!���� ���2�����'� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �B��[\ 3�1>2� �����������P�������    �����(���������"H����b��������(��"X�����������J D��� �    ����i������)�H/!�胺� �l��&�v���b���.uw���������     �  �  �  �  �  �  �  �  �  � ��� >P/S � ��&�L�(������2�������>�����0��7���(��t�����'������s����������8�@9�@:�@;�Jrr"rq"&�6(?���!.~ ����!.~ ����q ���!.�p �����q���o ����v���~��<�����n� � �&�d�?@��O��D1�� �*v�&�t�����"����t�����"����&�k ���)�����r���� .��r��%���� �      �����'��'.�u��o�ת�Ǫ��"��"��r��~�)�/��"������僜����&�!�������!>��  �P� ����P�e�O_be?g�J>d e1 � ~ ��&���f��b��BH��m�$H����"�����)��         ���jl��b
lb�j��)�l
�<(��H�H!���� EbFfG�H J�I��"��"��"�&�/��"���ߚ
"
����"b�������j
�k$����j���˪ ����� �&����>�
 ��� ����j��lbd
&!.��)��)�&�(�������!����
�|�J���(����/נ��h��������P��P��P��P��P��P��Z��"��"��"!N�
ǉ���J
k"d����j������������� �ں�>�?2��2� �������&�>�Pb� �/�� �>� ���Υ�f�(��֨�u��b�l��d�����/����������,� �       !��c��F��4��/�����J�����k    ���Ëh��!���i7ɤÃ�� � �"H��l�/ʀN�+ �"H��l�/րN�+ �"H��l�/�N�+�����OP?�P>� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �� �j�� �@����� m�m ��C�T _ @�� 8 ԄLMT_ ���3 ߇ �	%  � ��C� ��`1���� x  �  �� � XOReփ ��"������ P`�$��A �S��`F 	�Z2= ��Rq��C  �  �  ��w T�YCփ_ A5	�� ��"�I2_                                                                                                                                                                                                   �xذ       �                     �                   ��M���� 5� S� �                                 � @   � `� p  � �                            ���� ��������� �!~������>��ꪉ��
�b
�r

w

w
�r
�r
�r

w
�Y́�ɓ/�}�y1���?������

g

w
�|&f_f2[f\yi|e����f�23&_`&���w�|dcf^2B�v�u�'�I����J�/��"ӊl}��� �� ?�!��� 
.

������ u (��|u |%�� ���J;�fL<Bx�!`��� ���z�zib{�{-�������c�l�0�������đĀ��*P�=�Ā(���˴4��Pp�Pq�_r�Xs�W � ��}����tN&P�iL���cdb�d��c�������-�����r�|�(������,}��}j��t�c�%\Q@u�u@��� �� ����� � PI�5s ���)SfTJf�%b,iG�6I]b���{{�%!&�]����&��(��!!c�0�� �b 4f0@�0> 1:�1�    ba�"�S��!.SI"S]fI�/���J�k � ����&!"& 6" """c�!����!�9��/�BH�"�?s""��"��O�����J� �    ? ?`������ "��� �r0���]�/��!��&�9��/��r��zq"c�����������#�z��?���?���?�,�G�?���?�,�G�?�!�r��i������!��&�9��/���7������p"�i�I!r �&����&o�'��IT&�!���� $�� `/  n�� ���,G����� ��&��(�&�rn��g�"""br��n�!&!�9m�/�H����!�p!&!�9m�/�H���m�)��{ �!"���!"���!"""c���H̚"r �i2�/�!���/�غ!�"���!""&"�?�H��"�rx�i��p&(?���A�o �4i)3�&0YF�1^=� ��e ���&�^b���^�b�b�b�n��C ������{H����/���#�b�s��&�!�H����/���$�b�z   �&o�'���&o�*��*�&q�'��� �""��cs�/���&�؈��� � �	�"�k ""�9!���"��Hޛ�ދ 	A��Ћ  �A���$ ��	���� �8?f9@f�&��&(?2�/��"G�n��t5c(��7b67b66&6(?�H�!H�m� ��7"!6⠒�6�?��"��5����6565�/�?��.Ȁ�5!.4�i@ E�j7"!6⠒��8���/�5�4�i9 >4b�(/�������6�s5����4&�6s���� �  ���~  J B�3 D8 -�         ��⅂6��Bq(/�����C(��!4�����D���4�&��6��'��B(����d���4�'��G���6򅀶(?��66c(��H!���/����(/���(���(/���(���(/��l�"��+ ��&�&3333�J11b� �         ��� 0`������: ����� �]�/�"��!c"!w%&%!.!�/�"�c����,)"!7�"'G(?��O����S� � �]�HI�&]�HI .�@n��$��@�@�@�!��H����#lR&� �   �&/k��#r%�b�b�b'i� ��/�u�'$%&�&�&�&�&'כ �2�/�2����� �  ��	���оf��0�  & _�^�r n&r n&)�/���!1�1cw))&)&&.�j(����o�ê�����"�&!>11&>��!�s11&��p&�"cw>�_�������B������"c11&2r 2� �                      
 ��� ������ �__&^&B~i&~i~ib�~�~irnbrncrr11&.�j(����o�Ū˰����!>11&�?�m"s11&����cw��p&i"������"c!�1212b 2� ��P�o@/�j�� �                                    
�@�
 �		2�U2@/U�U1b؊��ȸ�O� ����e�/�2� 2��֖��6��62 .2�b�������ע ����/��"���!��r��ע��:��#��ss�Ⱥ��U�*K�M*)�Қ�Ҫ�ؘ �
�Ub� �    ��U"U�n��4(����i� �                         �GK���NJ� � �d�/����)�92�/vu"�Pr���t*)NSfXYfP�NM)NM&P!.Q�/�2����$/#&,G� ���
&P!.�nP.

4�JR�/�e��*)N�i�))S
'I
'J�/�I�����z�zi(��-iL��� �                                         $Wz!w�H4V�ά.��O*)KNb*�����ON&�))
'
'�N�*K�M*)���������P�"*N�zz��e�P�PNbOMbN~iM~i�~yk�X�Y����N�j ��&��4�c�F7�J� �                                                                  � �� � ���m �I�/�W��IbI!.W�&z� ��{~�(��~i-i��Y{.�{){)�����b��&��&�*9K�c*���ͪ��C��d��6��C��dh�"�hb��b��c�|��<��t��D��J�����"��b��&�!.W�/��������&��C��t��C��t��B!�����W&���                ��� Vf ��))
!>
c!�I!.(��bDW��l�<(O���,�<���D���Wp"bi&��tC�|�))Wp"
c�ǁ�
�<�|��K��� �����  �� ��������� � � � �� ��� �������b ��f�f ��b����������������� �   � ��qb�b��b����b�ǂ� ��o(��H����/�a����ư*��/�b�����!.��&�D�����������������    ��ob`�/��"

c(��
c(��
c�?����+H?!m����?��"b&�?�"��j   ��D�� �� �	^/I��2��b�c�!.1�/a� ����}j�`f"�����b��b�慠�}j��@.��ɉ����t��4(����|��ɀ��}i���"�����B!`�f�/���}k�����}���    �_�"����_�q���&2�/��"�l�'�B�|� �`���/��B@����`@C��@ � �3V4 �O�/�[�����\����OH/!��Ȁ��}�tO�@!�j���,}��}j�� �����&�
&��f��f��f��f�&��f��f��f
m2 ���/��!��!.��d�������/���b��d�
"
d�
��
&q�)������J��;                           ů	@ ����V��0 ���6��C�(O�i������&��5ҨO��ҧ��C�����&��t�.��b���.��c����(?�ԣ��?�գ!@���&��$�!���&������(?�ԣ����(?�ԣ�����sҀ{            �Q����P���������)��
�s
�y ��נ�I�/�z�zi�k�כ�w J�K� ��       r n�&�(?�@�!��&,�����8(/�����&��&>�*?(/�����&��&E�&��fk�&��/����Fʹ���&��/ك������4!��ʬ��!.��/���j ������"��b��b!�������!�������&�@/���          �V�| V�V�i� �V�LV�<� �!�� �@9  �2�/�u"��f��f��&��&���h���������)(����d�!.��/�Ǣ��b��crs��c��d͎J���H��F!�Ǽ(��b�Άǀ+ �β!�������&� �            �P�q�/�]�I)�S��]d��!S��~iI�j�))

4!
�!*���b@H��� � � R��ׁJ��� ���� !��c��F��4��/�����J�����k    �b"��?�!.�ba�#���&r (�� i�_�/��"��&r (�� i�_�/��"!�� �   �WǁW���� �WW&�WÁ�� Њ�}%���,���}i���,���}1��`�f.�����}k����}`��,+��}j���� �����c⨈��}�m����/�3����[/\�/�3� 3�fcD�����|�������c�l-��� ����f�/���}F��������2� 2�_F�&�������w�|���ފ������/�������QmbR�f�q�i�&���Q&����QlbR�k 14<�BE�MS���V<G�N\Y�P	rqD��[\fc�/�ڸ���[3b���c�/�ڸ���\3b���c�/�ڸ� ���㨛�X�/�Y����X�"��Y.��@��@/���PH�R�R�k ��W&� ����V�k V!W��������{ 	����Á��΋�wΛ ��d&�wÁ�����2!.3�/.y�|ڛ �B耤��+��� N���� ��f� �zz����� ��Pb��/�P�P�"i
&����
&� � I�]⠘�!{){)���� �I��0 �� `   ' � $��� � Q�� �� T 3�	耤�  ٳ� � �`��  � �a �N �  �( 	 0   � � 	���  @nL� �I @                     �                                                                                                                         !��bK�/�����K@/������K�H����/��D��� RD0  U @d AP�3�0K��  jl�5� �  X�`�`�J*��                                                 `����� �` � ������������ �  �             �             �             �             �            ��bf  �fb �   �  �  �  �  �  �  �  �  �  � `����� �` � ������������ �  �             �             �             �             �            ��bf  �fb �   �  �  �  �  �  �  �  �  �  �                                                      ���	 �
� ����  ``U``f��D��D                                                                                                ���`����� ��`�                                                                                                                                                                                                