���� A    �  <&	 << <19 	<7 <43 "=  -=  .<*  1  X p <���������                                                                                                                                                                                                                                                                                                              �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �  �� �� �� �� � �� ��  � �� �� �� �� �� ��  � � �� �� �� �� ��  � �� �� �� �� �� �� �� �� �� �  �� �� �� �� �� �� �  �� �� �� �� �� �� �� �� ԭ �� �� �� �� �  �� �� �� �� � �� ��  � �� �� �� �� �� �  �� �� �� �� �� �� ��  � �� �� �� �� �� � �� �� �� �� �� �� �� ��  � � �� �� �� � �� �� ��  � �� �� �� ɯ Ϡ �� �� �  �� �� �� �� � �� �� �� ��  � �� � �� � �� �� �� �� �  �� �� �� � �� �� �� �� � �� �� �� � �� �� �� �� �� �� �� �� �� � �� �� �� � �� �� �� �� �� �� � �� �  �� �  &��<� 1��	7� 4��"P -O �.*/ 1 ���b�n��&q.8/�H�&/&{�bb!���&&��a.�/��������a.�/��������&������j&&��/`i��bba���'��r���'�����n&����������66��J� �   ��ݟh�                                                                  �� �.�1�����.�������`@����� �o8?`�`@����0 �� i�b�@d�� ����N3�b�� ���3����������: JIՀ�Ѕ��0N ��J&����݅��0~b.����<}��بM����D��ب�f�����	������  b� r��r��y�/�����������������Ԛ��������������Ԫ|���|���J�/{�� ��	6ؠN�
6��C �d	
7 �Jؚ�F�� Hh  ���u��%��U2 8�J	eA�8��������&��z�z)!��&�)��yiF�.(-*&����*�J�썫���-&�Jx��,"d��� ��wiv".w�����uШx��Oxt��~�.�� ���ϸ��},��/���s��� �bc!� �J������!���&��� �@ BP����Ư�Y��}�B�������2.������-�ꭀ��(�r2����은｠�d�x��A��q�&�@.p/�@�o���Ϧ�s F���n bm�..b���B@��l&� �    F��k�&��� &�i�)�) �)��J� �� cb�J
�j F� &���؇��  �4�I����/���s����f����� �b	�l	(?� ����		D�	�(��	c�l���|��	� �l ���&�|� �J�/�|�$�J �,�h-�hi�xh�xg�xf�xκk ���K���bj(���������������i��
e ���������|A�d��ci��
��E PkbS ���b$� (V'&f�#�a���c��b�bdn0��bH(���(�����'��b���`)b����_i^�]Ғe��(�(&�&�&&D_Ӓ]Ӓ�&�e ������^_���+&���   �"bi
����(��#�j�'�]��b	�D(R]��b	�N&R]��b�W�Y�����9�3��܉و��(����@���'�(��!� (���������������/������ ��&� J
���� F� b\F �&�[)�`)�m"ȼ��/�!.f���bi�[)�b�	�� �   #���/�Z�pb#bDe�Yi�+6�|�3dK �!��C(���/����a���Э �H0� �� ��k�Xb������ WV)UV)��W�(U�(������|��K"�/�T��!�S"T R�Qb�k Rb�QbPb� b� �����b�Ob�����
�d�
Á(��V��N�������� �n���� ��������n��#����F�����J��/젮�Mb�L"�ք֠?���L�(� �   (��H�����f�&��bV���n}! ��	&	(?� ����	�J	 6  �! � K �����J�V)� bV �t���V��  Ni�{N��V�(���Ji ���V�����V��VN�������O���V���b  cV��&���j����d �  `�����)!.!�k|d�sظb�0�� �� �S����8f����@n����8@��h��(��I�H��(���(/���(����+��+��+��+�b@n�����������@�&�&����&@��&.�������J���&� ���.�k �!���N�6�CV��� t	c%� �)������  ������	�	&ɕ����	�z����	�j|r�dH����� ��� �e��	&G &�
&�	Á
� �J�	&ɗ��ƪ	�z� &�&�&7t D���	�j�	&��(?���(���(/��(����B(����B(����B�����!> �d���	�d	 t�㫮 ��Q�� ����c P�����X ��������H!� �d����d���	�dI0F��I0	' �J����&�}�   �����b �k|O�d��"�ջ���?�|��dK��& �,}�� ��̲��r"!f�� �" �l �<�����!�& �,}�� ��߻�|��{K%�����G��f��G+ԃ�idD�����#ai�%&�&^�%bcnH(��H(�H����� &�&3��� �J^�$�d���%&^�&�%"+%&���(��#�j���b	�b*�i� !	�R F��� F�!.	*t������G�4�8�M�C�C�C�C�	�	�	�	 p (��n ����� �����b�b$b��/���$���b�l������� & """Xo� �J
�
���i���!"!�c�.��r!$�$�b��&$�/�����b	Pb �l�݆�ކ�߆�� F��	'�� J
���	 t����� ?���� �      |��d����|i�a�c�� �khPoH��� � �iTbH � �!�!�G H � H.  &�� $&F��� ��#�a��%�b^i&%&E2 ��%\"^i$!.�/��&%D"+%&������C"^i������#�j&&%'&%D"+&E2���$!.&�/���'&er�ye"�i��C&^�&&&� ��a�i��k �Dbckw� �X�E��������%�cB�/�%�D+"%%b��/�|��dK%D"+ &  t '%A"+ &�%�c �~  &��b '⠡����z�!��&#D.ez)Bbb@����?-�*>b.�����*�JyD��J���ӛ��& �,}�� ��ܲ��r!�k � =  rRF��{�� ���t��it���IQ��(�<'z)�n!e"���!!.e�))bD��&T�S)2SQr�b�)rG�/�)�z!�b@(�-*&w�?�>.(�������*�J�y�D�!�)(/�!��|��dK'��&$�)'�"+&$!.& /���� ���n�k(/{M������n�;�/�٫                   ������������6��(�6��(�R J
� �bRJ ₄�   F����%D"		cE�/�%�	Zb	:y�%��&^�b�+"^i" %b	Zb	%r�& �)%�"+	&	�"+
&
	7
�"����	':���|���K����&���!��ؠN�6�O�<`��ث                �� � � ��l��6��?���� 6  ?Łl�(/��� �l��<�! �/��#H���J
 ��&�� F��b�F&�� F�b=R F� �j F� '� �|�\������"����V)��	�bcH��	�z�#�:ƛ�V)�ƛ��P.TI����ى�0'��  �0������ �?                  r��Z����66,6 �" ��|�� ����9%��9������k (����b�nbb��bwh�#�b#%6�!.#(?���%!>��/�%���J�w)S�&#!>��?������ᠮ#0����#�##s�%&�%'�!.%�"����b��f��&C&~�*� �� � S�F�W��� �� � -�	趤�  b�� �� ����  � �� �H �  �( 	 0   � � 	���  @�L�8� ����N � ���� � b�� J       �
� �   �"&�+ �04�9 �<A�FK�PU�X\�`e�jn�rw�|��� � �
���������� �   �������� � �� � �� � �� � �� �� �� � �� � �� � �� � �� �� �� �� �� � �� � ��F��� � � D�����                       �           �             � �� �� �� �� �� �� �� �� � ��  � � 0�� �� �� �� �� �� �� �� ٠ �� �� �� �� �� ������)��)��)���n&�d�� �� �� �� ̠ �� �� �� �� ө �� �� �� �� ٠ �� Ԡ �� �� ٍ �� �� �� Ҡ �� �� �� �� �� �� ԍ �� l'	�} '� ���u��'�xR�k�����  ��{�Ɗ��=6�h� ���Á�τ)� �� �&~')�J���s�@-�T���(�e�����7��D��J�����s���Ļrźy�R�pl"I�/���W��  %��U �%                                                                              