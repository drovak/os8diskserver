���  � � D    ------
--   3! -
	;	,";/* */*7+,
,-!-'0'	.";,
)%4!  ??)>���������                                                                                                                                                                                                                          b p2@ NDU_ �� �� �� �)�."9A!Sct�������hy ���sz�"T]"i�"L#� ɇCW;� 1�MN L#� U3m�%�H�A3� 0�SA�3"b��LB�1 �1�T@҃ � ��T@N� V�8L`!���� ��A��DUSA �P �� ԣ�V`�@�� DR(�� `PD0ăLiQ L�1 T2M��4� 0L#� �R@��F2E�$� �R@�Ne Lb�1 O3 � E�	5�8�3� Q���D�N� V�B3R�LB�1 �4 �S	�S �BR1��L#� �5TXOB�L2�1 �8�N�M�`L`!�8VCi L#� O	1��A3 Tǁ4`�3R�R`�3@�0 �NBT�	��ɇC8�MEN �TNT �8F�`� �B3R	�T5 �  �NBT�	��U3P#��MNQ LR�1 �0RC �TN(�d�OB�L2�1 S5`�""�	��XS�� 0L#� �R1T�	��XS�� 0�S�����	��XS�� 0	���C`� T�PS QN�Rנ3�#�4�E3 �BR1��L#� R���C	�S ���1 S�D@��� 0��3� �5T`!R���C �R �0�8Ք3	����;ăF@&� DS��R1`6�̓A�3� @� DS��R1`6ģFi& R �E�8�d�OB��3 U�NBTD`����L#� 	� QP8NR��C �BR1��L#� �`�	�S L�1 S5`�'���HA4D�m1UŴS�,X�8M T�8��CS���A�NB ER���CS���A�OA��T��	�T5 N�T�LD ��`�LD! P8L`!�R1��C��    _h" �      �8 �,(                                    ��x�1                                    q�R      �.1��            1� �;                                      ������0����ǉ���!��/�۔�����c(��Hr��*��c��� �������ۼJ��w�(?�F�����0����(?����� n��� ������6�(?�����c �����H  �
�����;���    O� D�0 �
X')��� X"'ӛ�?@@ �(�'�� c��� _���c��l��"��c�����r�f�n��k�&�6�6�6�5�����&Ȫ&����������   �����b�l��      ��/���͚��!.��&��,��� @���� ���b�����B�/��!����͂�����������d��K��i   ���7W)V��7�!�P�!�P�l���1���� >!��&�����������(���<�����9 �� �����������6��6����`_��D  VC``��D ���6��ǃ����{���8�S1���	 S��TO�#`7�@0 ��1�A�P@�AC@�b��2 U0�� �C �S�Q�1�1� 1�@��	/6 �� -,"ͤ��G*+ N  QS�&`��$� $O %� 4� �` � A� ��� C� C��D��D�`@�`@� C� D�`@�`@� CӠ4 %Q`0Q 3� CU`6`�`2� CS��4�`@  ׁ@�C`�`C�` Р4 ��� 0O 0O ��@ @��� �Ā ��  P��� ��@ 	�Ā 
�Ā  �Ā ���  �@ Ā Ā ��  �� @� � ���  ��� @��@ �   �  0!ŀ "ŀ $��  %��  &�� @@�@  A��  @B��  0CP�@  D��  @E��� F��  @G��� 0H�� PI�Č @J�Ĉ @K���  L��� M�� 0N���  X��� `Y��� @Z��� 0[��B  \��N ]��� @^���  _���  ����0����p��������������0����p��������������0����p��������������0����p�������������F0,���Fp,���F�,���F�,���F0-���Fp-���F�-���F�-���� 0��Ā ��Ā ��Ā  ��Ā ��Ĕ 0���� ��Ā h��� @i��N %j��C #k���@l�� %m��� @n�ѓ Eo��S %q���@1s�т @t�ѐ @u�� w��P                                                                                                                                                                                                   �  `�� �  h@0 � � �B P�V �L P�@�1 P�L@N5SDQ�R@�Q� 0�	 �QU�� �G ��@�4R�R@�R�  L�T `` D * � �j P PP��� X�E ��` ��$ Q��@��1L       ���ڙ���x�ph `X PH @8 0(     �	�������șǿ����������= �  A�4= �B�Ã= �PT�`O ŠT` ���T= 	���@�@6Ɠ1T= O�= À�  � 5Ã= �� �  υG�� H ��P5I� 1�  �  �=H  �
ׄ= ��.CÃ= ��@D S� @�#� �N�T�D � SƓ1T ��E ��L@ �TU= � D���`/ `
 �D  � � �R1= �D R� ��h� 1` � �D  �n.Q�� � փ�4�R@ �P��2�3 P�l ���� �� �� �� �� �� �� �� �� ߉ �� �� �  IwO�z w�xs js�I��p�� �� �� �� �� �� �� �� ȼ ��� �� �F
AA�AD�EV�@ 	 �1����D��E�OS@�4��D�FRX��    ����" �!��E  DU��#� 5�p:�� ��ENX�� �  �E�p
� � S@@��6 Ne@�T��C��0�� ��A�	  �������������������������stI�zw wO�x m��ވ�8�����
��Ɲ� DS@ �6��3 ��_U_�U�LULUUUUUS@�6��3��3��3��3 5كJ��һKTU�� ��0� B @���D�Q����3R@�P55O�1A@3 ���"  3//3��"��"ю"�"��"�Z#Z�2��"��"��"��"�\"����3��3��3��3Q�#��3��3��D 3 ���3��1� �C� 0��3��3��3��3��D 3��3 ���3��3��3�L0�C ���3�������N�@�Q� BP@A@E3 9D9<D<6D6DD99D<<D66D��D�@�� �� �� ��  � �� �� �� �� �� �� �� ��  lllfllfllfllfllfllfllfhif�������������������������Ϫ�Ǫ�Ǫȭ��� �� �  ��w��w�ֻ֨��� ��  ���̚��8�_����  � �� �� �� �  W[�RS�UJ�NF���  3@������	D��3��3�5��5;�[���޷��
�a�g'�n�'��DU�HD;DCBe��D�eAtN ���                  ���A      (�         ���A                                          ��	�A      .墼��      ��
B                  ��B�       ��oW                        ��� �   � �                            �                        � �        �� ���� �`s��������� ? ��   腀w,�$q�quUU��1� %w ���zE k���Pnxs�R�j� �;�jB�uo�wa���,�ż��B&l'Xie*�|&�&S:�(�
x��n��&�Jw��{	w��{	�'��x����u8�Z��ZZ�r���#��
��&k���Z�%ri��� �lƚ�l�P�:F :liO::�jS�~��h�f��I@�::&�9K 9Sc���Xf�7W	 �z���xޚ�p�� �x���� �p'��r��(�m)�a���X�g�{W�`�`�`�b�b�Wi(�����L�Z��f��h����b�b�iiY���V��y �*�lV���&dk(�� ���/��aU����a)�/��[�kiTX�τ� �����lB�/ފ�G�PB&���P�|��+ B���GB&���  ���F�&��&{a�h ����6XK 
�a��o���$��{�����dC��\i10fC�)/D���������0c1c���*�y �#�&��&� �o*�� � %fX1�K֨/I"I&f.�U��qʚ�֒H���[�v ��X���´���� �   nכw{	X��
b�H.b�&kՖ��K�{���&�#&"&� ��������9=ll������ˋ���/���B�j�U��X�&zK������&Aj)   �
�?&�����6��#�KcK�/�<��i�`)V��� .�`)[��!`�W(��!._U��cW�.����)[� b��ਁ@��A&?'f(b��������� �	�&�&��4�ji     {��\�'e��7E�| ��4��GU��?`)X*�&zKn��w;�{	UJ��U��=��U��;�!��U�<�*U��f7��U��f�.�
U��.�".fi+(���U\��U��f�1�
U��f4��U��"��&kT��U��$���*U���"�U��>�~bIb�jW ��JX[����k`��J�U�/WY(A�aV���
U(�� �
�KY	��@U鼸�������Ui��UϘ�X�U���&k�k��)`)V���)D.FJ`)�J (/���W� ��X�[������U��U�kY��U���k���U�#X�U*�k(���X[�[�a[�k��)C `[��[��Ě�*�U@�X��Xi�"���a)U��kT�� �XU����ki���� ��d�"�B��/� 4&zKn��&{IwH�0{	n��w��{	��+�jn��w��{	���jp�=�jp�!;�n��w���{��ju2��u�5�
n��w��	{	��$�p�<&�p�&&�g���(/�/z|�SiR��x��n�������z �)�/�f�.W	�]��1�Q.f+�� ���4]� k	`���� �� �᧞��Ib��&n��&{Iw��{	��&�p�= !��q��=�/���  ��q��`�X瘗 �)5b/6b07b12b�3b�4bƧk�)��u�/�
2�&uD��n���k      f$�/�/��bf���f�A��&���i1&0&���y�� �v����y� ��<� �OP^� � �;�Sg���B��K��@�HW�
zȿ{{������&n��&�Kw���o�}b�j�J~	&>&D�8!�D���}&&1�&0�&/�&&&����J~	&>&qۚ������J��Ib�iq��`v��JX����[��X�� ��1&�0&�/&&&� ��	����    �	;�SgGD	Df'�p���@i��� �
(zk�{�{n����&�J�w)�{"��&k��o��c��0c1c|b%fef�.W	�S�R���x����w�	{	��Jz � q	{��(�kw#���st����m)v�Ƽ��/���<m)v�Լ����m)v�޼� ��� s	E"���� �V��� �W ������[�l�%"�o�>~b	dC�	ǁ��JzD��Db�/� �����(���1.����{%�%HN����.�.�n%bF�bCl	m.�%�J�/������m)v���� N %�Jlm��/���c%��%�mv� N�%�� �])])])V��])Z!���/�٫ ���Fp��G���K ��t�'�&��@�<fU \	$(/����;��/�,�h�$��;�1Q �.&l��� �,!.��/�(��@���� �,�&,�&(,b��@������ �1C D0�� �8/&90&:1&q{�� ���4c`�KW	��`ś t	N c%�w�s	w��N%%siw���
�&�%�$� �`[�l�� �!_�[l�b[�l]�����F�.��$�������?b,���c����J.K�!0⠱�1F q��0�����G (X�G�"ȱ��!.�/��������G (X���(�J (/����j��ɉ��c�c?,&�<��b(��CF��O�!.�H����b!�����/ .��b��/����,,&��J� �    d	H,�,�k#"�@ f 3F � ��� �� ����� �� �� �� �� ���b�L�Z��H!���� ���� � �O�� � ���f���?�����j���Y����?���Y��    D�/�s�� ����%�J� �ׇ�%O�[�� ��n1 %�bQ��.Ⓣl.C0d
��cC�J
�� �1�K@0��K 0oP/"/�k�s� ���H� ��l�<�H�N ���� ���bd����(� �N(���@G�V��� �(�c�
F�
Á(ϻq���/�
���6��ã�l���� � &f�b�bti���h��ဎ������J{I�b�j�&� �sw�$�N � ��c��x7�K F�� �J
�
�� ��O ���F��4��h��wS�^w�   /��,�|�è�V������l�<^��&ʝ��Vi���V��X	�V��X	|&!.�/�s�^��V��� �!.|�/��K �\���O�(���(/�ʴ�@/���@����"� ���,�||&&st�E"���� �V��� �C�� ��� ��� ��&��r��� � �x `	[��� �����������������l�����W`�lO��lyP�1F �`9�l���
l��(��P������_�lc���lH�P(ې������y���D��M���i�l����� ���y����������lY���l���	� �   �Y7	.9��Y�R =�S�g�� `	[�������hͮ�ͮ�ͮ���l�������&������� �bh����?����������؅��� �D�湹D��� �� ���� ���4̽c��F��Á]�̮DĽ�   l���͋   ��&��Á(��!�l�������*�� �� �lR��(/����/��K��E�S�  �P����pP��Y �l��(��C&�������(�����U�lO�����U��lyK�	���W�����W0�l���V����w�Q�l��w`�l	K������ྸ䮸��D��&������/��l�KY	�l��������/�������7������[)���U闢l�������;����C &���x @���=����� ��Q J�aV���d��U	QVY��K�`��a)� �   ��4c\y���!�K �������!�k ���H� �Q(�&�w)N.��D"���� ������������!I"(��@�����ހԾ*@  �l��O�(��H /����� ��������*Vi�y*FkN����� �F����� ��� �gt�sw��#�����&�!.��/{��f���f����&���?{�����j�N�c���N���*��(� ���&� ��{��+ }f����t�w"��{��}��ks���si�֨s�� t��bK' .'���k d	NZ	lN�Z� ��<�k��jP P�� f����w�>��{��{ � bI�/b!�Ȯ�"����"�b���i�i��bii�j�ߚh)h)h)&�ߚwB�	�	��bb�j��Á��&�*&�*�l��<��1�0b�/�f���{�h)�h)�{�i��i����� �I�/��K���������� � ����� ��|�K �&�Á�� ��/��K �st��	& �l	�< (O�!��/�����K @"n"�k ���� � b� � .b �&� ����w�%�{s��*� �t������g�{����&�k �/,&����/�`U�_XI� �            je�V��X� ����.b��J.��������"�n"�.�j ���h���{�B&��H/�P��j��!�@n.b��O���.�j �/���b�@n�+ a� .A�d� �a.b �A��K ���$/�n� ��.ǁ�� �.�<� � � n	���&�+��&kiw0��
�/������*���� �kE����� �lR�F� �lJ�K� ���bD�� ���4]���I����= �lK�cW�*�� ���<P��	�(���z��ÁK�!��J�0J
��!.�!>��s�HT�����  ���F�'��'�ù���e{E����F���������l��|P�'����K�FÁ��(��AAbj����@&F&k�k�k�k��/�����s����7�7��?�����r��|�P0n����(��n�����!;�����0���(/�&$���&�&X��/��(/�&�&��ŷ�n��$ � �/�?�!54U� ���� � J��J�����b��b�
c(��
c(���ǁ��Ç���b�hs�D�/������Z	����� b�(/˫����E�/�&��/ˊ� t��  J\���{�  � U� � \
� ��  ]  �h � L�R� �� ��\��� ��   �������Ӡ����Ġ���������ƽ��8�