���  L �E7  ���������                                                                                                                                                                                                                                                                                                                                                                         ���@�bA�bq�b)�b+�c�+��&�&�&�&���@i������� ��b��{ ��á�d�
>

����鍊� ��(��H���)귛 ���6��B���@ �q   ����}��'`�2c� q	@љqК@��Ϥ@�qϛ8!4Р@@�?�^]��NDO�@� �������BIF_&t)�) �q)�q�@+��q���@�1���&�&��&��     ����b��&��Á����?�@�7�����
�l�
'�
'�
����������� �Ψ/�q�@���̚��K��k � ���/�!��� ���/���ڴ����� /�l�q��}O�HH0 ���u �u�!� �X��Q� 	 4�
�����@�␢���r��c�����"��j   �����/�@�E+���l��[�W���ݼ�� �	�����{ ���4(���@i q	�q�@q�q@�������@i�q�� �! f(?���"@����!�/�@��˛ D.  bDD�  &�  !$� ���K��j  �P�OD �d8y  qJ@  �	����)��)��)��)��)��q�@�����@������!�����ǁq�)0�)J�)W�)j���à����'@����@���������s���Ƞ�� ��q�)�)9�)P�)C�)[�@���ډ�������ǁ��@n�������@yv������ʉ���@y������������1	K�QO�Ofx���q@�������@F��������q���)����q���è���&@:�q����?�@�P���?��"�@i����q���è���<� & �6@��@ �@�����������9� ��)�)�ؾ�|�2�J&c�bbb�j!.�/�b��� �Gi�F	�E��i��\Y�:� ������FDW�@ϔ@'����q@��������!>�q�@���Ù���q���Y� ���������b��b�o�@n��"������⨲���&��"@�����D�ˢ����)�ò��������     )u�)�������&�� (�����)�����)��q���'q�� ""
.

�"���nwPH�Y�w��Hτ�Y� �t �	��ǁ���ğ@���������ǁ@ɝq�)��)��)��)��)������!���ǁ@���������ǁ@������������w��� ��!��&��?M�>L�=K� q	@������qI� ��� J�� & �; ������D� ��)�)�)�/����ߛ��p�i�!IH�GF�EK�QO��Dyf� 
��6��L
�t���� � �	��(�q�)��)�)#�);�@���� �bc(��� ǁ ��J�&���/��"D�P�����<�)�M)�g@�F�������ǁ����?�)��������)y�)�������)��)����������'� �
 m2�V�dHY��N�DK��?���@Q�>f� ���)�)��)ɚ)ɮ)��@�{����bИj��(��(��(����� ���s��¨����D�@����ǁ�� �����)�����7�������3��|�� @�� 	� ��� �   ���&� �� ��!6׉L �< � !D�׫ ���7���J���[ID ��PfQ��� ����y !�b

c(���/�@�@	7
��&D.�"�@iXq�@1����� ����� f�b$�n%#f�2(���/"6"�"(���@.��/���"P.�/�#���/�#�H$� "b����  7#�J%�J$�B�#����� ��!��&������k	6���  ? ���?���R��`�OXN�? ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �          ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    �������    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����������� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �          ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����������� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �          ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    �������    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����� �    ����������� �                                                                                                                                                                                                   