����  �C �  !< 
8!';
9?>(*%8';% : ';?7> 
 
';?6> : 54?3>(982?1> ;(8';;?';;?> 

0:?';	/? : .;/>(+ 

< 
>(-,+*/).y): )*3?<!>% > ! !??                                                                                                                                                                                                �������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ ~�
��D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �� �  �����}���v	P�n�_��Fn n�&J.
�����ȳ��������R.�i���b!�⨫�Ȁ����}�� $0����&W ��&�@�|"���J"��&���|����/�C��J��B(���}Ɉ � ���k   ?��������������������������������HB�?������� �/ �� R�` VV�!�ڠ/�F����ڶ��r��x|b�i�(��m�������(��m(/�@��|��i�����m(/��������z�� �"�b� �F.��+�(/���H��bV�������m /���ڨ/��� ����� ��c�(�������F�� ���-�����?8��W��2d�pD�F�&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{ �(?��B6� � �gWq���� g�t��D����/���}�� $����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ���������  @��    �bH�
��bmF��B@���Pn�����彀�O��O��������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�׷�����2X��(?�
�

��������������o��R1��D��� N E��D� �@C� ����	��T P�ل�MA	O���� 0���/a� �&�	&�	��J�g�v ��V���T� � � �? ����  �;> +':'9;'9;%'8'9;&'8'9;''8'9;"('8':$?.!'7.!$?.!6%'5/%	  	    :   :   :   : ????????{56<683 8!3 8/4 27A: 0 ?=<,/,)#�������������������������������6��6���H ��� >Р�����c�c��{0(����bm�/mm"��bm�&��B�f��Ɉ ����k�c�� �������r`���O�֮��&���Γj �   w�?���&��&���?r��/�V��/����yN� PT0B# �텿��f����dw��DW�b��f�Dd#pD����&��) ���"�����)�J��� �	�����������{�
��*������/��"b��

d
(?��
1�����)
�9�������t�����������+�P���)�h� ���֣ � � ��  �/���/��?�˟�!��.�F$�@R��HH�V� �ɇ��`���o��W�>�����0�����S����0�����) ��������"������������y���E������B �A�B ��I��0�����������Ø�E��(?��c������9��`>�?�/������vÀ�� ��KW�x���P�O���Z x@1�Ywh�`��'����` 솀�����R��c(������ ��������+�����b���!�⠺��2�&�	&�&	7D�������7��� �� ��l)��  0��� ������ � ��@?ڀ��"�b!�@��d�É���Dܯ�����J��� ��=����c�/?�� �ɇhY����0�1������8� B�B��A�L���  0�L�	��@�L��� P�L�
�DC �vE�	�C0�vE�	�B1�vE� ����1 ��V���A �vE� � �	ct�᫣�z�����?[���#H��ϑ����Z����� 
 ��c�g��w��7� �����!>@/�
�� ?��
�J�
� /�	�
	&� ���É� ��� �������"��� ���c�����/ﵛ ��&��������Ɉ ��c�/Հ��/���k��dS�������	 ���{���F8��;��oyO;`\���썓D��D3̒�D3̒�D3�3�3�3�3�3�3�3�3�3�3�3�3�3��n��&��'��0�����)�ӳ��P(p ��b��&�J.����b�ۖ����J.P����U����"��b��&؉<�@.�/�����&��É�Ơ�� ��b���� ��ے�����)�����; �         �?����{ ����ů����� �KNUk�U������P��	�Ф� 8  ����� @3������ 0   !-6{|7z"7 �z�#�/g$�t� �u#    �� �      �}Ɉ 7	�7<��O�   � A�8� ����������������?���� ��!������ 3����� ���@� d�s���������������3-v �l�&�&���@~�����&7�㐋��	� ƫ ��  �����|�/�//D//D/�N�}Ɉ .�ؾ鐈!�l}�� ) ����|ɡ�b��hP��!��}�A /�
!�,ˀ�� BH��{�rz�~�y����z�xP�Փ���l��<� ���&�yÉ
Θ���}�   �
邼}I�  ����,�- /�w�|(_v*�w(��*�X�*ubtb"c!*⨡�"�J�/vs��"�rq)w|�p(�"(?o$��n�n�&!'&!,2���w�Po�m���hÂl}@���lt�$$bp ��X.��/!�x!����"k0�!'$�J'j;P"F�i�h�+Ii(g�**bf"&*e"!*bd(&!�;�ӛT�	݄ě���;��<� @������%!.cq9|&R!q�|o[  �%�&-bp(�b)�w$��
(᠐�(�?������)k F��!.(/�!�&���a4>X��8+�`&� ��?࠮&_&&$'&'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[�   ������i� �;`.       ���/  `  ��ˀ�� ��� �� ժ �
 ����8��������	������!�#%�')�+-�/1�35�79�;=�?A�CE�GI�KM�OQ�SU�WY�������                  PW�Z_�bḛ  ��������/�%`�0? |/������m�ih�������X&�k��%�&��Ji�h�����l�lk)�%���d����h�������mY�lk)�%���d�h���������   �����	��ŠTP P�!�s��&sK�*!��"��*p'+o',�+ ���f�h���n �bD�.Hs�b �J��)�� 4+&�!�����c�� �����)�!������#�a"bb�j�a&#b&�����|_&�\6�'�d\cc`&�`�a�/�`�b`&���jh��`�k_���d�J\�Jc�Njh���ik��h���jǚ������ժ��t����s�c�*���/�-��b�p�   �
�@.b/�F�u��<82�� �瞙 ����wc�"�@_�����%@����'���>�#��'��9��2��s�����'��9�N�����s�jy�+�h+�i)kh���j��+j��,�h,�i)kh���j��,��>j)�-�h-��k9j��.h�.��kj��/�h/��k9�N�j��0h�0�ik�h��j��0���u��2λ��Z�0�	/�	�=�
�d�<;"NB �TE �TɄ�8NA 	5I�3 �T� 0� E��HMN"��T� 0�נ3T�8�`I�3 P3  O> -\ K: )     NB �TE S(�D	AcS  � 	���4�DI�3�[��C�/�B�6I��&69����B��X��JB6)b6���A&(?�6�����������b��b��b��iV�9 �	d�9�j��1�h1�i)kh���j��1��|_&j��2h�2��k_��j��3�h3�i)kh���j��3j��4�h4�i)kh���jÚ4����'��7��� ��3�j��5h�5�ik�h��j��5�����D��� �9���� 0 ���=�(�#���Z-� 穞�� �Ʌ�D U �C҃`�4T� ��q	ȃ2�mKmm�mm�mm�mm�mm�mm�mm�mm�m � �	�$	�3�L Q�   N� S�`C`Q�4N�`  m�mm�mm�mm�mm�mm�mm�mm�mm�m �� E T�8�`3�TB�� 8 N��S  � 	A�� �
��)��&�@���E��� 0�H>������d|b_�b��k���b\ji�6�h6�\k)_�J�|�_ji�7�h7�i)kh���j��7d����������b\�j ��a8 !V&r�B��> ���@�  �n@� �� ��  �.@�1@�1��1 ���d��6� � x �ۢ�݂��d͊���  �������J� ��w)  J
�
�� �H� ��	������di���#��"�a�j���`|b_ji�8�h8�`k)`�N`�"a�/���`_d�j��9�h9�i)kh���j��9��a�"!_�`ji�:�h:�`k)_�O�`�`�"����`&����&��&�`��!(?��й�Z
@ �� j	�;�h;�i)kh���j�;d�������t�$�`��  � ��	������c&bd�b\�n|_&\���\& `&j��<h�<`�ik�_�JdO�j��=�h=�i)kh���j��=�����\b`�j��Dj��>h�>�ik�h��j��>��&�d|b_cd������qp	  rp
  sp �^��D���^p���^q�� �X� ��	�(����c�n|_&�&�d_b�!.]]d��j��?h�?�k��� �`ji�@�h@�`k)_O�d��j��A�hA�i)kh���j��A��j��Bh�B�ik�h��j��B�c�O�c������`|b_df�������	�  ^s��  �������H
H����䰙
(���
7�<��X� �� ��������\�n������d&|_&\`&j��Ch�C`�k��_.__b@�����`�d�Jj��Dh�D�ik�h��j��D��\�!��(���(/������\�J���`�j���\�j���\�j����N D   �N�DJ@ ����C  R ��p] 5      �h6!   �� �0 �	������
�b��n|_&
�6j��Eh�E��!��k_��j��F�hF�i)kh���j��F�����������. ` ������������������� �/�8�N`!NB�T�T 	�R1�D��� 0 �bc&�b&].^]&].^.^]b\���+                        ��fʯ�� ��	��������#�a"bb�j�a&�b&���\�bc�n|_&�'�d\b`ji�G�hG�`k)_O�`�dO���`a"���`b"`�jj��Hh�H�ik�h��j��H�cOр�\)"\\b��/�\��\&��������*      
  ��`�e�Z�J��������T P           �@�� ��  ,�	��������#�"�cb`�n|_&j��Ih�I`�k_����j��Jh�J�ik�h��j��J�`cD��������������#�a"bb�bc�j�a&#b&�c&�d�d�N``d�`�c\&\a"���b\"\ji�K�hK�\k)�`�'�/�d���/�j��L�hL�i)kh���j�L�� ����_�
�  ,	�	�c�ccb��/��������)�c&�c�_'bd_b``b�H/�����!��\\b`ji�M�hM�`k)�_�__b���dO�`����\`&'d&�j��O�hO�i)kh���j��O��cc&c(/�����������V��ʺ                                        � @��� �	.�xB��c���`cbd'b]cb!��__b����j�P�hP�k)]�J�'�]�n__&_�/���j��Qh�Q`�k`�]�J�'�]'b``&�d�ddb���j��Rh�R�ik�h��j��R�c�N�c"��������X. �  ���� ��� ��������� ������%��� ������1��� ����<������{��? ������c�n|_&j��Sh�S �k_��j��T�hT�i)kh���j��Tc��ʨ��� ���|�_iikj��U�hU���k����_��j��V�hV�i)kh���j��V���� 	���ʴ����AG�8G "F��@R�N�!�T1�C�. �QF�u�7� �P(/i �O�� ���<� ��	   � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ����H.�e&�"��c�n�g&��?   h	������=z 
  8 � K� ���(��bJJ�J�茀k  �   ��b���F.D����"� �    ��	6	 ?��������&�{  ����&��b

�
{��[�����[�� � �	� � �j��Wh�W͒k��� � m	����&��&� ���b����"��+ &!�����   �����"����pݧ�W> nb�@  [0�� �̃����Y � ��&�!�ʋ �"��ͷ�� ��L���� ��:�f�)����?�e�)����F�g�)�������������T�  �R���C� � ��	� 85<N�`N%�E� @〮�P"PPb�H/���m�〮r)� � 5  ?� Q��PSɲNB��穞 ������������� ���b$H/����!�z�&�(/�z�FF�F�⟆k��*        �	����j��������j����������j��������j�������j������������dǓ�Z4�#�P����FiBښF�BޚC� �d���3Z�J�������n�ջ�� �� ��� �=�� ���� ���� ���� ���� ���� ���� ���� ���(� ������� ���(� ���(� ������ ���� ��� ��� ���LԲ������D@`Ra��D��; �� ���� �� ����                   穆��� � 
 	    � ;� ENB�TXA��	�3��[�D@`�c ��HҠ3D��DT� ���H�`C�Ʌ.R �H��C	��R��KNT"A #A�3LS ��2   ������� �������� ����������� ����������� �������� ����h��� �        ��U��Q�ɞ� ff�)��0��c

�
��'b��biikj��N�hN�i9kh���j��N������ ��� �� �� �� Ϯ ��    �� ����ݴ�ݷ �̷�Ѹbعbۺb�b�b�k��⾿j ���� �� ���� ���� ���� �� ����N%�PE �S�  � 5�N ��`1�/��%?���� �� �������������������������K ����� .��d��J��d� �    	B1 �� H �� ��/�� �������'��; ���6��C�(�@��

�
����0(���@/��"�۔� �   ����� ���&��'�`��R1�� �D��@�?����� /�! � �� �����;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    3<}�tq�on�m{�| � ]�cD�HO�i����g�ܛ�ۖ��y��{�ۢ�������d������� � � ��������� >��y������ � � 0ܠη����@!�������� ���������6��H��h� �   ���������; �� ����������������TRN�!   �����Ⲡ����I�������ʘ�6��&�ʘF.���d�ߪ !�/����/����/�������������k   �BR1  � HP������ L��!�� ���� �