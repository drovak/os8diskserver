����   B    8     8
     #  5(8 3-  		2  		 7   <<   =    <(   <   =
 
 (
    9$   <      <.                                                                                                                                                                                                 y 0                                       6^ c� ��  ��p�" ��   ��)#    o t;�	@ @  H E  J � 0� O� F�T��6  Y��Fa   P  S @�h  �mA  !r�F  �w  �|� 0@�A   ��L 0��O�3� p�Z3���   ��`�  F��� �` �`��F �CME  �B��    ���� 0����@� pRa��7�    �̐D  �D  � � D M �D  � � D 
�D � �DM �D � ���@ 
 �	�P �`	�� 	�MQ a	�� XT
  E#E��@  @0�  !@M &@0� +U 0 0�U 3� 5U M1 :�U 3� ?U0 D�U3� IUM1 N�U3� S��
X� 4
  ]��
@bSEJg�0kl�Clq	� jv�	�Ci{	�@o���Dn� Pm���@@ ��@�  ���@@M ��@� ��Հ@ ����  �AՀ@M  ���  @ 0�C  ��,H���KƁ�GFˎ�@UЁ���$8Ր�0Gځ�L�/ߒFL䁓�T�R�%X1���  ��� 0��  �B� @F��$�`  @ڀFF @  	 "C  
 L  	 8 "Q 	 %�! 	 *"� 	0/# 	 4" 0	(9P#  �>�P 0F�CP#�` H�P�6F MS#  �R�S 0F�WS#�` \�S�6F a�# 	  f"� @	Pk�$ 	 X   ` u�   z @�$   �� @�S   ��� @ �S"�Q �S%� 8 �   ���L ��$  � p� @�L   ��R  �!  ���PA�Q�B"  ���F  ��F#  ��� P   
��   �C! P��rC8��T!�	 H�"T 	@��"  ��A 0@�3  (� 04  H��T
5�JA(�T�5  P$� `  �  .�D  �3D0 F�83D� =D0�Fa B3�  "GX1 PL� 0&Q4  $VÁ3D [�44@ `��5D 
e�46@ jÁ7D  �  ! � P  � ��2j�        AN2  ���2�i�ߒ����2����ߒ�����8�(�(�(�*�٘��8ߨ/�F>ȕ��ݠ/�����bgww���(/��(���(/��(���/���������7�����K�'� �G� ������N�/���� -�p�����/�	%��!��k#Y <�����0͎� ��	�2�             ���=� �                                      � �        � �                 b{�  � �   �  �                     ����a�P��_@m�M� �!�dh?P��`��* U��UP3��K ��2�/.�/1�/���6&~6����}��|G�4�/�4�D�3����a&{6&2�i�(/���(��(����6t�����/�|�2 a�3b!3��&1�&&a&/�/�}����(��z�/y��HIF�J楠�//&�J����(/�J��/��Ȫ�&13dĂ�1�j����4D��Qs���v�� �? 8�6&@�����@.78b8�7.6�J78b� ��!.˞b��b��k  ���̠/����O����F.����7�J.
�����r��d��J��)�Ŋ��&��BɁ|� �   � �   F&�	&�6&�Á	�6�J� ����z���c��ˁC �            G�@�����$�� ��� ���&&Kxi�}���� ��w��H���!⠛�!>�/�|�D�;6Rr�|��� ��*9&+:&,;&)<&}Κv�/yu��9�*:b+;b,<b)wi�H����''6�0 6'�t�|��t��(��sr	,}i�v�����q)���c&�l ���"U"&R"�\"E6"0M$�h�3t�� ����T ��b&fu����pt� o���n|���=��"�(?�('��#@.��/�Ϫ���� �'�/�|�X�+���$n &�+�"�/�#�@����|��&p)t�"�/�#�@�����#��m�&p)t���$�n&��
���$o ���|��'�/n &p)%p)t ���q%�#n!.$"&��� � �e��.&����n&pt� u	|������ ���h= b��>?&'b$b%}i����y�'�B(�h(�H� �q.&�!⠸�@.o�/|��� ��6&�6�l����66Co666G���66&a.6�/���� �"o �X��՛��t־�
&��
r
t{ {Fki���N�� � ��W\�(7��  �|�T�� 2���2aB�f���(/����EI�J�j��EI�n ���� ����E��EJ����J.b�1��� /E����ic�H�)I�/���EI��I��E)�E)�J&� � ��dĀ6�CЀ��ī ��i)���Ћ s (���H/hj"E؛ &!����������&� ���F��(I��������D�0�� �w f� �!�>�n-�ix��wܚH(��6���>Co"�������Jy!����-(/�H�(�/��H����Ϛ}��� /��"b�"��: ���m,�(/{��6�0�>�"6#6�!�-�"� `� �4D; D''D=�/�6���6 v�!�|S��	&-}i�7�-	C(��7�/-�j��_}R��@ �	"o ���@.#&"�"�o!(����n#q.&"�!n�� �k" n# �"� �"n #b �#&���#!.b�J�"�#b���a.#/�"��"�*|����bxi���q���/���� .&&}i�v�������&&O�u��ܺM�� �@R"����#�� )��(?��*a.�?�+�a㠞�,a.g0����B66cl�����: �� ���K7'*'+','&6&w@.m�/�f�� @��f"#f�蚀"b7#b8�h�5����@8�##&7�""&݀�o���H#@.�#&"�"o��J��/�"Bo(��/�|���; #D#�"."o��K�\� �&���k ���K�������j��4���� ����kv2 ��(���(/���(����+ *+,fѷ������/����)���H�*��*�*�h�+��+�+�h�,�ʈ� ��ܸ���� ��ڊ�P.�0/р���K ����@������K�܋ F�� �

�
s����
�F�%0�]�����Q '����-�h�&&&n F�&�"&�kUS�VQ�Z`�_ � ���6.�h !�{� ��.�`�ȹ��~)�~9�~).�/�~���D�D� �(��f��̜�����(���~�� ���(���?���J���(/����̷�333333333  �E)鰰  Xn�h �������� 3m ��Kf$
.
e�(��$.b���M�n�$��'�'%'�ɘ�t�LKDɡ(%�(t ��.b ��M�/������rMMe�'���1�/��n ��dj�EɒdK����~K��ɘ� ��K������N�/ڊ�N	�gN&���/�4Ob1�nHIf�J��bXnf5fDLf.�K���ɔb� ��(���� Q �9�.������'G�/���.�/���.����cE&���Ji�@�  ���� &m�{ !�{�|��e &p)t���fyO .� /�(/���Ⱦ�f����K#b� ���/�#�DD�%b#%D ��#&|E��#�b�#&##6#f��|��*C_�/��|i�b�c�� �k�h�PH������Qg <���� L�-�&-�i5&5�I �5�bH-�-�#/!�� �	���	�b�b6c	6t�{�P6�� F�!6��rw�D¨������N�      ����Mf���@ P �`��O� ���a �
.
e��6&6�26�ln 76cn!7H/隷��66t�6�6a>�/��6�~���
$����������)��I ��/�f�d.�/���7&�Á7�7m"7)b7�{x��w��H��o0���|E��t���x��w��J��|S�t��nⷁ��&x)�wϚ!���� ����6g06'6BF�6�|������66������o ��ob.b�t�M�n��

�e�rn'�t��t�� 򀈒Lp��O1&t��5tk}t�!7�t�r6����6p)�6�pt� ��)6)7"����)Bs����n (��/ ./�l}��v(/������y�� /u|C�/�k!�/�������ઠ�/xi�q����/�j�/��#&�ݚ����#$�`/�!�p"�"�䉬#���!7�18&p1�7�J81&t���/\Q�_�� �  ��&Ԡ�ԃk ����ԸJӠ/���@������z
�
�⡁l� �  ������&�� D�� ԏb��b�j��O�b���Ə���c�J
��

���J�0��d��0�(/�����ˏ����߉lҁ<(���N�  b����0 z�Z
���dҁ<��d��k         �;��������f�� F�F&�FÛ�i��/��ߚ&�&��,N� b��,N�� �b���y��K��[ ��(/��B��brz���&�P.��/b��� �  �b�� �.�/��������z�����/�c)c���h�s�!�����2(���(�FÁN�� b� � N����N�mN�k꠹��D ��K����[:���LM ��/����/����z���  }���(/- Oh��y��``"&�b�-�����f����i�� �� .��*}���(/���H���|����J���(��@@�1����b�����XX��Z����_-b�����)7�a7�7�7d��p9&�Jt ��&�&t��Qf
_-
 ��R� C�\�_S:� S�R&R!.Y(/�����(������ ��7�77C7��J� ��C&��(C�777�7�7�nCC&�J� �Z�/�Z�Z�����7�7�7�7d���YY&� ���(Z�/�7�YY&�	&��&�&��d�7�7t7	7�J��(�������Ë 7�&@��          �����Rl
�_PXY ��y3                                                                                                                                                                                                                                                                                                                                                                                             �8��'''�r�b
b!7��6&�&	6
(?�r);�l	<6�<�i;�<rs6�l�<�l	=6	>6�8���<�H�����<�H(������=n (>����&�6&76�J�"������ww7�J8�J�6&6t�������n0(�����w�{!Q&��3���:�#8 �������N���G�@�� ����{P0(���"&"�?����Ĝ�����{{r�b�r�rw��ˁ�ˉ����O�L��G���,�������N��!�ƾ���s�~��y렞�QrN�i����(?��'�"6�&�	��#&	7#�J����{�ö���39�8y7�  ��ESݎ�D�D������'��'��'"b(���J��H���J�&�	&�) ��	'"� ��c	s	v"n �c�J
���"H���J�&�"	r��	�{�`�D0 � � ��3 Q��S �QS;CU�T JNFBMRAMKYJNJ[LA[GS[PO�N�D;C  pF����  �hiQ:��� hg� � ������6���z��(/�����㰰&��<�����'��'��'��'��'����'��'��'��'��'�&��K      �����&��/��������"h �
�{P0�"&"�<�/�|� ?ى���0�����'���!  ��'������*��1���yp���0c	�8邁����A��� a���D�)�����"H�����q�OL�)�m����6&)�n&)b7�l7(?�7�7&&�J�&&)�(��~��~9��~��6g ~�z�c~��n0���d9~��)�L6�J��E���Ʊ�������������������ж�������������������Ʊ������������<y��B#p��� |D�5