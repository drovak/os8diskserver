����  @.     :09=80*27>(*2$*'6$+8 !'6.!  $*>$+.4$1>
=.4      > +
0&0!+0"+6661+62: .?    g6$ )	)
)
0 ?<h   00
=	; 
 ?>(**>> *%$/$,(3$,(;$.$,(>8 @ S@���A �3�< �0A @ � 8p �<,� (,@$$�  <�$�?�$0C,
 $ 3�  �$�?�<,�?<A/� < 0>� 34,�?<��6C ��2�*$@<�4<@ ;�3��� > �iy �;`.:" � ���/                     �   ��w��w 2�;��D.������� ��a� �������������������@ ���� �e8�@6�� #��W���`��/J�"�
�F��! �?��A����2�  ��������/�%`�,D�-&��6���$���$���$��$��$���$��$���? $�K�, ��$���$����8�/$䒌 Π$����$���< $����$���: $����$���; $����$���7 $����$���= $����$�����$���$�%���&���$���$��$���������ʄ������A���������A�/���� Π����A�/�%����&��̛��������Ϣ�������A $���D�/$���$����$%�&��̽���������������A $���D�/$%�&�����ڬ�$���$��A�/$������������$��D $��A $�%&�̼����������������$ɜA $���F�/$����G�/$@�A $�%&�̼�����$ɠ�F�/$� $���E�/$����$����$%�&�����Ȭ�$����$��A�/$@�L,������ڌ������ବ$�I�/$@���$�E�/$��$�����$����$%�& � ��́����$����$��A�/$���ϐ�����$�@�F�/$��$����$��$����$%�&�L,�� � �������$�I�/$����$��$�����$��$�%&�̼�����$�F $��A $������ ��$�E $����$���l�� ���$�H�?�/$��?�/$�$ ����$ɪ̔ ���$���E<"�$��< $��$I���̔ ���$���H8"�$��8 $��$I���̔ ���$���E7"�$��7 $��$I���̔ ���$���H="�$��= $��$I���̔ ���$���E:"�$��: $��$I�߸�(�u� !��&��<�� c���̔ ���$���H;"�$��; $��$I���̔ ���$�E $����$���$�̠$�%&�̼�����$�F $�����汊�|�F�$�� $��� $�$I�$I����扲�|�^�$�����/$����/$�$ޔ$��A�� �
��)��&�@���E������������暡�|���$�����/$����/$�$��$���n��l���ɣ?$��� $��� $�$I�$I�格橒�|���$�����/$����/$�$��$���nՙl�����?$��� $��� $�$I�$I�����  �������J� ��w)  J ��������������栊湂�|�
�$�����/$����/$�$��$����恺�|�$�$�����/$��?�/$�$��$I���恂�|�>�$���E�/$���$�O$��$�K�,J .�$��$���$�%&��́������䬬$��A�/$���yÉ
Θ���}�   �
邼}I���M����栈����$��@ $�$I�$I�$ɠ栜����$��� $�$I�$I�栮����$��� $�$I�$I�$ɠ������$��� $�$I�$I�$��������$��� $�$I�$I�$ɠ������$��> $�$I�$I�$�����;�� ��������栈����$��� $�$I�$I�$ɠ栜����$����$�$��O$����$%�&��̱����$��A�/$���Ό< ��$��$ɜB $����<�/$��$��$ɜB $��,���8�/��$��$��C�/$���8 $� � ��$��$��C�/$�� 0[�   �jPU��$��,���?�/��$��@�/$��$���? $����$��$��@ $��$���$���$��̫$����$�����$%�&���ʴ���̽����$��A�/$�� �����������$��> $��$������$��$����$�%��!�.!!.&�/�!�&�n*&M,6"%&!!. ?`&���DbJ� J
��&�/��������$���F�/$��bb�&!.H/𠯠(�& .F��&.�l$���&��!�$�,$yJ.�!��/$��$���o�!��/$�$9�!��/$�!�$��O���&�J��̈$�%��ˀ� �L����c &��̅����$��F $�f�"b!������&�&J.�bȦ&�����<!��$��D�J�n��&�$��!�$�!.�/$��$�����Ɣ��� ����$%�&6�"!f�y�$x�$��z�$��$�'$�!�/$%��"�&�#!f�'$�!�/$#���_̈$�!�/$%�&�#!f�'$�!�/$#��^��$�_��$!��$�%&��#�!l'�$!��$�#�J^_̈$��]�$�!�/$'�$!�$!�]��!�$�^_̈$�%&��#�!l'�$!��$�#�J�]��!�$�'�$!��$�^%�&���]� $��^���$��_ ���$%�(��Ұ�����������ǁ  ���f_�Ȁ�K    �����&�C�� & � �� &!�k � ��2))�� �� �)��� �n�Bl��AϞ4���6�/ɔ��$����$� � "��_����"�/�$�!�$y�$�x�$��!�b�  ��������� �������ïظ����������Ġ���� � �� ���)�����������/,�+��./�)���3���K ����� .��d��J��d� �   �
!�A  �� H �4 ��/�򲮹������'��; ���6��C�(�@��

�
1���0(���@/��"1ߔ� �   ����� ���&��'�⻵����Š�������@�?���� ���� �����;��A����b��c(����?�����J��?���1��1/���K��C�����'��"��c��k� �����}�tq�on�m{�| ����Ȉ�Ԉ� ����������y�����g/��Ӏ��ᒠ������d*��+��� � � ��������� >�{����Ž`҉g���@� ���IJ� H��������6�-I��h� � ��1)�19������������; �� ���,)�*��+�����TN"�  �� ����/��,i�.)�1)�0Y����b�0i��F��6��J� �!������2�����2�����0��{�1)/��/疮 � �` �Š���ο HP���� �� �HJ�I��ހ F����&�� �1)�.�撆J� �   ���1�� ���1)��J�� ��|�A�|�����*��+� ����� *	�+I�1���b�ð 	��b����&,!��"��Ѷ-��ڲ�޿ð �� `� >��b�8p� ?��"�����'��J������ ��.��pݧ�W> n �IJ�H���� � �l�Ao��n��&� �����?�/�,3�,;��.),>��.),A��.),D��.)/)�ȱ�3��)ȟ�����y����
��A  ��LD!  ��N C�� �Q�> �����   C!�T@��σl8�$N�! R��D�	8�T5V�Cm!�PB	�C@R���D�8TT Q��PSɲNB� S`Q�` �@0	�
(@ 9�<    �<� 8 <	 0� +@$   0/   ,�+(�$� �4@$,B0030�  
B#,�,�+6��    C �0 �8
� ,  `0� `<< @/8�6�? S4 +�7#08�  .B8$	`.� �=�0�2��.4