���  � � � ��+"3*3.6+.	*$**1, *+**1,,,3  ,  -" 1)$	 >  4 4 0  "   ++& 		 	 	 	     		 	 	 	     	           	                                                                                                                                                                                                                �tg 
�\ u   �
�w  b�C��s b��'�  �twg ` s   \   ��w� p���w�7 �u  ����/w�? �����w�? �g ` �t �hwg ` S
SV�\S�
" s 
z* s 
  ��נ p�b���w� p�bԝ�w� p���� ����� ��b��
B� @b�Dw�4 ��b��wC��O �� ���� b�7��? bi�Gi @bfD�ft bn�gn `blD�lt bq�gq `�̪�Ҫ�ت�۪������������
� �z 0�/ ���� 𓇪� ��� �
� �����/ �
l�� l
�z���� z ww�O���w$ l
��� ���z��� ��z�p�� z ��/ p
�/ wwpJw$ �
*,��/�2Ǻ5,��:�;�@A��E�G�JP� ���� ��� �
� �����/ l
�z���� l
��� ��z�p�� p
z 0�/ wwpJz 0w$ nqs�vy�|n��������������������� �� ������O �
� ��� �
� ������O l
� �l��z��� �ww4l�w @l����O �z��� ��z�p�� p
���� �ww4p�w @����˻����Ի������� ������O 
� ���� ����� �l��z��� �l����O �
zp�� �pw�w�O�wD w�p*ww4
�"�wD ���� #�$)�+,�/.�48�7:���� �����/ �
� ��� �
� ��� l
� �l��z��� �� �l<� p
�z���� p
� �p�� K RVX�    R[X�    ^`a�    dcf� ��� ���� ��R� �
 l
< �p�� K                                 nq�s �                              �̪� �                              �������������������
�����������������y����"��$������%�����'����� ���� ��z��u� ��z��u� ���� ����� ���� ��u�� ������� ���� ��w���O
�$� ����� ����z��u�� �� ������q 449�= �66ݘ6� ��z�   �z�� ��0�       J      L��� �WW�Z\�WY�Y\�^Y���� �
 �� �C*+/��"J(�
���6��X����� ������3���T�K C��i�$`R� Eه��[sQ = "��+�PI R C D    I R C D    � � �       	                                   	                             �b�� 	 ��    �                                               ��    �               ���E� �      ����� ���!� ���`�s� 1�k��� `�`� � �@� W�q�B�FBJԀ6+:������� ��jf?�� �r��r���¨���� ��b��b��b� �פb��b��j ���§�c��D�r�� @ׁ<(����b

�
����r���(������ ��Eb��bFb��Fr)��J� ���b

�
���(��� �� �G)� ��G)�G)� �����HII�Hx����@K�*I��n? �� ���}���� /M���l�<kVE�V�y�L7�yH!����yLi���y�P�yMib��/�y�D�⭁n� �J�VEAZi���L�� �
 � ۾d�ت�ۢF�����rJ
�����7�&��D�۸����d��'� ��(/���>i� � �
��E��&��&���� 0 ��� �@a�h가�� ����`� ������>��� ������&��&��4���E�/    �'�''4���'�''c� � (/�F�r"�N�� O	����/P"��6���(���Qi D��K f&&666R"����I��K &!�ʀ�����(x���/�ٶ��f�θ@�@�@� �X �X@@������  ��� ��L� � �� � �B P ��dn� ��"��c����'��C��� ��E"(����Q�y�������� S	wU9�� �a.�/��d���M�'�L�<Vra��I�*&W�M�M͚�R@ PKM�Z���Mib@��J�T ��,\]���D倫�p� Z^bȫ��� R&&666666R"���R"Ȁ�����/�����&�)&Q+��&� ��"����/��b��Qi&���k ���F�D.��&���(���d�<��6��è���B����/��C�Qi �(?'�s A����WT��W���8�J �X  \�M12 "�/ ��&��4�f�Á(ϴH����S ��Á(ϝH���^�_]������U��U��
PH/����ob�b�j� /�Ţ�k������
[��y�J   ½����Z���E ,@��Q �M!��h�JIZ��I� T	�My�\�]ޛ `	�f��/�����QW��W�ց�� P�G   B�� ��d@>�/�����(���/���(���&��a����^���0(��b�ڰ�1!.�/���c)]��C�ld_)N)���_Қ�!&C�l.ca�������c�+r)!r)]����"�h�*��\�⨉�� �r^��øQ �S�lk �@� �' �(3 ��1�/�O6$e���Vn66�^��(+r)!r)]��^i�_)���6^��6�������_),r)D.N)]�� �cf�r��g�g"&�(s�� V E /����K ���&� ���@�� �"."�d�ʫ �t�KX� @�D� �� 0�L� �@���R � @���tAu�sMH�I4����4Tiq)Bh]�)�NX�/�*��h�I�T��N)+r)Fr)]I� -(��zZ�$Xi-�k $^���_I�k�L�� ��/IQ�I�y`i����/�����QW�M��"���)-&y!.P�()h))]IJy��M��\�]I�W	� D��&T �䍱L P�V �C  �T��ԨP 0%٣����k�*pi�Ԩ�t)''D])�z)�$XiIp��f��/f���W�X@����M�.�l�<VR*"b*c�d�66T>R"�����&Q �S�UT�To��h)]*�Ik ���FV��fn�?��(��w�/���l�<b��S�
U) .�Syw.4��&U ����3��EKM �((bD(�&&( N66'.�lZ���i)c(�,���D#F��'&�l�_�#�#F.F��cH���&��#&&���c�l(2���(�&
&D�D��C!
㠩��(����d��f���&��2����!>�?����#��'V��n�I{    H)� �<�o:=f&F.F��ߠn��tf��(r �Oi�/��&f�bcdn�?��b��G�/�S� U	(�&�����'B�yQ#��I�WӔ B����<�(�a�?�kZS��L�<�n&U��T��&rFr)]&��'I � �r��� �R �P 6� � ɉ`) �;2�'1
�- ��bb(b(��d.cd6@>�/�����(���5&�5Á��(��a������D�C�(��zC�& �T���<c]�(�/�T��jrr,�r�(d.N]�& ?�V�&z9Q0���S��U�D(�J��QiBT�w)2h]�)')tQ#�� �h+�r��L�!r2>���Ok�Z�?�/�S�
U)Q	T�w)2)CFCh)]Q�#��Ál�Ami �IT�
#�c�]Q���Z5ၨ���ig�55cׁlT�d_)�N)]���!&T��!r)]�i��g&����<.r�|.'.7D� ��br��r�Nכ $^���_I^��q2�   A�/�A�Ss�]� ���P3 ǣ ��g���S�@�Sk���� ̘�#L�T @` 6�W� ���1�K� �	 e�� �@�@�@� �R �R@�B ���B@P� S	�BlP��&U�Q�T��La0��� �cך�d�_���<N]��Q�kI�M �Ti�jrr,�rd� .�^�MN�]��I� ��e��
  �n� �U� 8 ��"��&KM�Z֞� �I�4b���4^I)h)�_)]��tb nIkM!�IkM!�Mit�JIt�d��!���TIqCb�Lc ��lClf��&Zၨ�؁��?� �i)�!>�l,rr�!"�o9s]�B(^i���r�NI(�J]�a␭��J�W���@��z��2�/����Qia.��h/��u�~�"h����k�n7(/�!�76b�l6�<�&Tq��_),r)T.N)]T��r�c�]7����r�������e�:  ��F.�� E"�lrrb�|u)uG�rbN��rviQ�� ��c�_I+r)Tq�jr),r)D.N)]�U:!]m��[� �k�x�b6c	c�s ���76�'�7163626D62����	�		b��/�	�������f����,c(����?���b���s����'�V2���� ��Y��.�����r��ǁ��� �a0����� r�{�u)vx�慵A�[�ͷ����� H�S2P�@sadm���������q�vT)�,�r��1c)�,�r1�]��������߀������ـqt�3�(���l3!>(f٨���(�J�3�a(�3&R"(���o�٨���O�(������������&٠�Ӊ��0(tʁ����� ������d���Z� �٠Nc)+r)�Ál� ����iq @�{�|V�� ��ݮ�������)�_)+r)�0�a��.�b��/�d��1�c�������l(?��&�''f��Á(ϼ�� ���b"����������)��J���� ���^��_]������s�(���S��]��&(?�!�c����J(?��ց����G��q���ۀ��D 5� n�?- ?����� �2�/���̀ހ�y߀��ܝ���������3(/���3�!(��l(�"����
����w�7���Ca����T��N)�_)]Q�������w���xT
� �c�]����(�JQ#�2�/ډ�1V0��&��6Q ��������g� ^	�N)]��w�=� ��Ál���"�Qi ������O ��N��P���^e�N]��ܝ���߀�3(/��������w�7�w��3!>(�l���6��>Zn�� �i)�4�O���lT�d_)N)]���|Tw�� �c)](����/�Q����2����1�01�r�������Á�������Á����D��J���:� ^iN)]�j�������܎��a0������w�7������KQ#�3(/���3�!���(����bi��!>(�d��D�<��b�(b!���j��&S�U��(�J�L�<lP���(���tTywd2_���N)]��z 0�g� T	v ��,c]��\� ���������&��Á�Ȱ �    �t � �S �U��� ��8�3�
P,=�˪>� �(����������� V1!.�E2�j�r)�r)�J�װ u	u�u�u�uv�� �e0���&6���cp���cا��0t6��b��ce�'�C�sr�w�|�U�� �e0����N6�� �����'C�.�{    �λ����Ż��D� ���`ꐐ� ��q�Ԫ�� Ъ��Ī�� Юɍ� �D�/���wqD��s �2(/�ȿ���q$���q��� ���j ��_I+r)^���_I��?�^��_9�]I�Ŵ�  �T� ���H�K0 � �X�K00 ��S�k� �� 0�E � PV �Sl@����ˀ,�@��@�@̘�n 1 ��  ; � �����@.��/U�@�Zᨍ�6i)�&�6'6�L�T��r�]���t�B�{Ǩ���1!.�/�2������"��lT1��,c]�� �e0�����d6�T�q�L	6	c),r)�	��f�r���(]���)�b�lg�g"&�<os������@�>_�`4�n���   ��l��&��&�c)+r)Tq�� @��<lg�g"&  `Z�ᨫ���4e������c�漁<o��jr),r)s]�� ��0�������� ��d�6��C��F��(��bbr	�b�l^���<N]��J��	�r!��j��ˣ �� @  �0�������T� � M�3    �`�� ���d�&�&�"�l(?����i�:D���� ��2����T������c]��L(?��&(?�!�c����J����R�� �3(/���3�!(���6Z���VN6"6B���l)��"o ��"��(�ȿ����  �����/���    �fV���n�`�                                                                                                                                                                                                