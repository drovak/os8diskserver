�X����&<��̺��[:���׎N��x��w2m�նN�S䮎�F���dRE�2Ԯ�L�9G�E���"s82dh.Ɨ6�n�&'�&���D�6>t�4�e�1��|�"�hۛ�kދ���rBV�ðqc����dΑ���d�A8� �<^��b~@�Xe��zgꢫ���3�����g[J����@�U                                                                                                                                                                                                 8   �B��A�^F���  0��F�	��@�^F�	�  @�^F��� P�~F��8 0�^F��� 0�^F���F �^F������^F���σD�^F�	�1 L�^F�C�	 D�^F����^F�D�T  �^F���T�^F����^F���P 0�^F�P�C  �^F����  �^F����^F��T ^���PP�^F��� R�^F���  �^F�S� �^F��L !�^Fߋ�M���J���1��E��T��E�U�T  ��D����֕L�U���@�-E�����@�^F���� 4�^F��� 1�^F��� P�^F��   �^F��ӀL�^F��ӏL�^F����L�^F������ ����� ����   �	�@ �^F��� 0�^F��D  �^F�� P�^F�D�r \�5C�� P�vF�����2օL� ����4��F�����@F^�����@�^F�����@�^�����@F^V����@D�^���BB�^F\���@ �^F� ����� ����� ���� ���� ��������� ���������������������������������������������������������������� �  � ��N�ԱD��N�ԲD���D ���˄ ���D�������˄ ���D����C�����������C�����������8����5����� �8�eߋ�����5 ����4 �����M����� ���������TA��L�G�#�������������	����9��������7�����P ����@ ������@�FW���S��FG��8 ��FGΆ�8�N������ ����� ���� ���� ������,.(���� �       ���'��l��� �����6o��������/��������/��������������������P p���!�扮½�c��d��6��B��b��l�?��s�!�Ǩ?��� ���D������>"��j$Г�Q���$Փ�$��q2 ��i`bgid�i����g�J��J,�����iB;�*����@�� �q ��"����l6�m6��6�l�B&h6C��lʄ�Q��Ũ�$'l���x����-Y�$'����-��m�*-�-h�����/�()-K�(��+,��j�h�/�Ũ��� � �i*)-ś ����ʻ�C��#� ��8�L5`I�C � `B�T@`��X����� @o�� ݦS1Iw��0pm lR�H����·�.6sX�<��2b��i����ٍ���r�����Ȅ�$딦+),���  i�Li�,����B2h�cn�co�c�߸��
�s v�!9�F���̘�6�6��3 ^

d����6o̣� F� �� �|� �����c�o����|� �$w� '�s @b�h�y�)��p@on ln�D H����Y0��s
����"��y�A0��~��y�A0��&q .��b����Ӛ�E0pqbD�!p⨮�p>"4p&�?2 �c�op�  r� &pE ��bH
���& �0� 'p�&�X� ��� &p� �r>�&��J��Ā �� �s�� b� �q .if`g&�㸏E X
l ����n�op ��@��U  �    q  ��	&4�&��	�r>�& �J��&��&ߘ���	ǘ>"��d�ߨ>�&�	����>"��b!�⠲�4�&��J��D�q� ���	&��&��!	� ��>"��b!����4�&��J� �����b�@n?��׉�� �q .��b	4b� �                       ��?n�P�� �f�b���ccbG���6 6cE 4�& �̉l�� �(/��������������� ��/��cb��b  ��b�k�� ����= ��&�̲�Y����= ��&�̲EH
����k � ,�?(O�)_� Pb�i������Y �K()�E0H
�)-�� �.\�5[� bÅ?kF)f�� �a=�`K��  .˽�˩�����������˪��������������������ȾjcD.E�4�&b�bƽc�����cb��b  ��� �  Dbn�cb��c�h �O�쐴�c.�b�� ͸� �cD.E�4�&�-��-Ǡ �?��<e�4d� ���;�"�!i�F������;0H���o ���'�7�	�t��p��U uT�%�R	$)H�4m?uTRe�-,d ��>�mu�U�$S�R
 "�H�mu�WM$ҞR1*�R�mu�W%՞Rh��\g?3��WN#��Ofy?�I��q[c�݀�/pm?u����zm?uS�ME�$"/sͤA�p��/�z ���mu�W&�b	&.�f�寺 ����mu�Y�$Y�bf廵}�9P.y9�H��m? ZM�F�
" �/�y?�I��q[c�݀�/�m?u������g?3��WS#��/�m?uS�M�D�5"������mu�TM$�R4�)�1���mu�U�%��R+i6� ����y��I�Հ���	�;33C`3t�J��U��� n
�i����
b���h����
���|���g�JO`�gib;i&�P�z'��DNKw �sO������\O�$�p�}�9�R���/.gO3��WQ#��/8tOp@��B��P�� ��b�����f����b5�}�8\��j��zd�%�����qM�e��1�|v5�m�
���izf�}�8\��i��b�"��u����u���e��)�xx���z�fd�%�����t���}�X\�&�ܭo������� xs�e�� ���"��f��i�O� ���"`��/����D.��bH�����$����"����b�����+       ��!��?������&�&�&�&��?�/�.��bЊl�
�@ ���'���	  �/���/���/��?��          U
{�<���	�������	�� f�b�n��f���(���/���" ��(����/���嚀����"����H.&/���t���������&������"����?���h�����h׀���h�����)���9���� ����)ـ�� ��Kꀞ�+� ��]�=蛮��S �뿾�?���A�]�� ��/����/��b�c(��(��������︻����6��&��9   �
Cݤ�@����F����������D� �  !�(?�����D��� ���?��?�˻���W���b��"���@�(����i�=����c�/?�� ��QT ��� Jq���� �O�V�x �&�(���p.oN�� .�{���@�����P.�/��K�����&�&t����ǈ�(/���(���(/����Ǹ�����(���(������<�����&�����F���|�"(���kX#
�, ��#�� �.��qߧ�W� �`��� կ
F� ���6���"���¨�� � 
.

����� � (���� ��(� ��(�(�(�/�������� �����o��)��"����.��k��"����,�(/��������*!��&����&� ���c��F��É�ȁ�É�����뢨��� �   ��(��(뀸� ���}] Q��� ? �I� &�������6��)� �����)�������cb�����)�)�)� �	D�� �	L�� �	T��N7��7PR7 �4 �T��D �D 7      ���l�ˊ��(?�����������Ѻ�2 ���J��+ ���r��{         ,�}V�v�` �� U*q��!J����od Z �	�� � ��/�������ŀ�  ������ �	� �� ��6��'��)�&� ���4(����� ��b ����É�� .�/��� ���(���(/�����ǉ����  �����i����� �  �������  루��  ������  �	 �   7�/Dq������� � ��X̎3�K �	�����涃l� ����H���b��i��/������.����@N��,� �� n��&�����0��d��0J
�
.
�� �    ��C���P�`�V`V�`�Li!�`�`@��k�M� �������ҋ ��|���ỉ��ʀ��&����3���� � ��?��q�T ��'�����  `         ���� ����� ���c�� �� �����e �줈��  �¨������ �$H����+,��� ���ǉ����;���18   �q� ���&qD.
��
"t�
"@�����������$���������{ ��V1x̀�_�O���y�����-�<-�~ ;�� �b i-�� b�$�����qb ��i`bgidi�,�����i*)-��,�g�J��J��˃i�;�*M`�d��4�ʂ!���@n��"�����)� ā ����� �   ��'��'���6���b��y�c�b��{|�0 �      ���[� H0 �/���) ��Yo ǩ ���� ���    ����(���(/���Ё���|�6�����6�(������b�����!�������ÉΘ���F.������|�<�(��H�����!>��<����[���e���]���n�� b�$@����&��(����)��+ ���ǉ��a@ȿ0��:��U�[�8��3�P��  �] ���� � �(����bF�����b��&��É���� ��b��&�J.����b�ۖ����J.P����U����"��b��&؉<�@.�/�����&��É�Ơ�� ��b���� ��ے�����)�����; �         �?���� �         � �KNUk�U������P���� ���?�������FN���&��,��|��C����������i�����i��������(�����G �&��� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d������ ����� ���� � (����B���ǉ�� ��������9���������>���������ɀ 5���K(����� 5����� ���s!� ���)��)��F������< ������~�f�i�/��́���3���&��J�*���G �偼�|�Y��`�ˌF��:�?߇( �UN�<1��?  ��/�����b��b��g�'Ӝ'�����y�&�|���xE��r��'�>�����?�����FӨ?��0�����0��s(���tƠ?��������������� �	���(������<H����)��+ ��bg�J������|؞� �-�������0� ?@�-�v������k��ߗ��                                                                                                                                                                                                 �;��V�            ��  6�	$��2��"��$ �o���f��f,�t �D �v��f��frdJ'uIG�6�  4N   	    8 ?@ �� �� �� �� �  �J`HP`��������������   � �� �� �            ���   } � � �t 0�� ����	�yr�k� ��� ��$�����$��!�F���^$�����$ϑ!��F��b�$ؑ"��qnqD.q .tqb� ���s�����'��'��'��'�ʚ��'  � ��$���ʚ���w�$����ઠ����r��r߀���w� ��� ��� u  �P1Q���s���f�O� NRT��$ˑԀ����$i��������$yg�������$yj�������� �����'��'��'� .Ϡ�����r��r��rҨ�����r��r��rҠ�����r��rϠ/����r�,y� �        	'\�2]� ^��D��������������? @�� �6�>�L3TR38�3A���3%3�?� > �	6	
6	 6 �0 '
�J��Kq�(��!濝& &�	& ?  s�!� �?��� �	�JO���>�&�S�� ~ �⑸k `��'�)����C��#��V�SO"�#1��A  �������O�X� ES0:w@���-?N x������
�s v��8��O?`��؇��  ^��/�#@�À^%L��qb ��4�&�l�_
&��)l&�
&��)�l&`
&��)���!4⠯���D���>"��j����O���� � �(��>� 9���=Di�i�"���l& 
�i4"�i�]�/���l n
ib4�)`�&iiB�隠i�
��V`�
pb���ܶ�o�"
mb��@W���@ �|�BL���c��� �(/������ �             �
���������(/������ �             �
�Ū���Ś�(/΂�Κ� �             �
�ߪ���ߚ�(/났�� �             �
����ރ��䳑���z�������xwf��x���f�ndl��� ��	&	�6�eb!��Ș��!.xf"Ȗ����/f�&'��	 �o 	�	c���	�	d	�6�G��{�&|�������EҠbD�E4Ӡb�����R����d�bf�b�����lH
���;�"
 n��&��
�r

w���x� ����d���         ��rxb(g�h��}�g~bh�j&(�2�?2���B,���� ��������bn�c���(���c��lH
��ƟD.E4�:b�5��c&���rw� ����dD.H�E4�db:5��c��&!�Q)���cr rbr�v �t�A�!��"y����Xa2xry�/��&��y2c�2��/���c�b��  �rb$i��L$�� 7�4.OA5O@-O�~O#qO+no-{O* @ $Y� I'�� o$ޔ�$�u�ng�nh�k'Řn�&o�zVnp�&z� z�'И� �p�&lB"zoz�?Ż ��&z /�Ũn�&o.zoz�6z_"zpbEH.
�zzt�z'zzGzpb�lbA�&z/��t�z0����� p ���� � 6�� @o!ii�%i�=��(/`���iE ��bH
�!q����4"j�b��&�l6��"kjb�okm6�m���� �mD.E4nmb:5��c�o&o?"�nb�o ��p�l� � ���y����"� x��?� p%� � s�� @o�k �퀳� �i�l�&���j�魯����� ����U�e��U�lUI1w    �Ӹ U�T�@�	H��2ă���>��� @��@   x�/�w�!�⠵��!Σ�/���a+�<��l��惠�x�l��bw�c�Ʀ�l4�&�V΍�'�����/�$��Z$�$�wY ��h��<*$��R$�t��'����$��RH
�)$� �RA&��+��l$$�wY  �H+)$��w��i+9,P���h,_���f��?�ˤĄB��̤���̄oC�����Vnw&��!��hw&��?���������$͕�+),�xl�D�2�� �  Sz ` �C\���� �(?���O�&,�-^���b(��(M�(�+����J,�������      ��&�
U�� y�r�b�g��w��~��~��~��~�Hr��b��l��fxf&2�&r�$&���Ѐ���$�s"i���!.q�/�D�4�&#�z-i�z��+� s�vOI `Lzd���#��%��z'�-�K()�E H
�)z�+���'�p�&#�Yl"z,i� ��� �$ݔ�� � ���ِ�r��"�/    �� `��d� ����D�فh�ٲ��K ��F���h�Ⲕ�K �����X�H-'-v2 ����^(/�a����,��-(9��4(��@��-�?�$���6$�;��亀�-U2@��>H/�ê = L()� ���b
�ԉ��ً ��
.

�ٔ��-�� ��J�(�� ��I()��J� ��K�(K�(�� ��4�l.�?� �!�à����&,��!�㨊��4£�l�è���/�� �yd f �����C

�
��ɺ8ɱJ F (��Z(/�:�HG�K()�,�� � ���݁ls�Jts&3u&uuCH���u�u_��a�"��j J�����b=��D.��&�
.
:��3"ʁl�`0�����r��r�s��{��'��'� ���r3b�r��{ �q�/>�"��b�r�r��ǁ��q�/�벍�b��	Hb	'�	"�r	'	>"	�d��������&��&� �      � �������&��~ɠn��~��i��'����M�Rm�( 8:�� �I�&y7O�|���'e�\G��U �6����    ��@�.��                                 �v'   SR   Έ  0                              �.(� P�D ӂK� 0�[�ͻ                                                                                                                                                                                                                                                                         ��/�$���$��Orρl��6�:2��i���E����y�H���xL���#�����#��!���x"�����-!�� ��j*,��()�-I�n�oP "����6��C�Y�[_�OR�^i�oq�iŐY�ˑ�.X���[,]���Z,��� �[]̀��\��Z��� ��^,]���L�� �]����� ����8_��w��w ���4 	�� @  ��˂��� � �(���j�*��&$���������b������R�/���H��b����i��b�����'�Q �������)�������'��&�����/�����b��~��)�����������b�!R�/����r�b� � �          �� � a����������   �b!����>=���& �
�������Ҫ����!�/������!>�/���������!�����6� >�?������c!����/�����!�����6� >�?�����!���� ���!���� ���n��&��'��'� �    ����������buj����9�( �	����b���Ҁ+ ���$
� �&��� ����a.Ӑ/��K ���6���� ���cѬh��K ��!.�H/�q�֐/��N� ��ʂιk ���&پ���K�΄�ص ��� �         ~ �	���ߡ� ���홅J���'������Hs�|���EGq�]e�ۨ�ջoϠA�Sjt�j �cLqWFs�=|Kr�h�
�Q�om?� �����2؅
~�K�z�RN1���A��lc�H�0��e6m��b��e��a����"�J-����G	:���	/��?�����#쀇���u��j&*v`�K��%�h2 9k�~+lꦙ�~���]CQ�u��ڣ��/ܰ�y/�����z�23͈o��kj2���,$� )>��0� o%$���*$� )0�;o� ������m&�j��nb��b��ɠi�
���a��i�������7�Қ����b�����(��t�������� ����d������j�&�
&���֪
�J��z��3!��� � � ��� Yl�+ �Љ��@���� �A?ݹ�D �  ��& o�
c�ט�9��b�ט�/�e����(���4"�Vnn/��s��y
�6
�<��n

&^&O��H ���������װ�o>"
jb��i= @�&(?����9�ܘ  ���J� ��
���� ��4��l��6��C��d������|܊���� 怼�� ��"��/�l���� �(�6�� ������V��o"��i0��'�zĄp��¨������h z�p��¨�u�����h z�p����il'l?"
jb

r:
&m
'm�+ (���pF��6$ ���K ��b+N�(-� s�� �۠�#Ӛ��jz6� ���6��)���   ��K 	��
�� ����\�� �����k�y�(ώ��4�&Vn���S�'��ő�� ���i��b��/��� ����/���YH/��������龽b��&��"��bF�����b����D� �       UpHb�p�ƀ���k ���(�y�� ���b

�
X������bF�	��&� ��Pnl�(Y�lc@��lD�
�遬������������"�������c��c���	 D B �AD0RD  �P ��'��'$՞����q������'��'��0Q�'��'�$���阶���$��������'��7��'�$�����7��7��7��@�b� 0�# U �� �MA���5����5BR1 �BR �;�6� �������̉�T����$������q������'��'��0Q�'��'��7�$�	���������s��s�$y��顫���'��'�$�����r��r��r��{ ���r��r�{��&º� ���s!������D ���« ����/������/����J�ް�%��(�2)":�s9� ��8 &CS���37rF�,������O��T�$��$��$��$�����                     AN2�8DkQB D� ���X(C� S�R��D`���AŠ��c  ��DO�#�8(�#S�`C��E`V��� �N$ �U`���� �� @�΃�CA��S�E.1  �B2���T� E�`P��;Ʉ�8L`!�� ��P� �?$ ���48N�PӄMDQ� �                                                         �d j j d�                                                             ������������`���������`�                                                                                                                                                                                                