����  � 82$':&��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                               �4�5������� ���L �       B �@8                     H �                   (�0��9/�������ˡU� � �?���� ?� ����@��p � À0� �� ���� �0��?�� �� �� ���������UP  ( 08 �'��ڪ������f�n&f�$�('&����/���Ĳ� ���~�&��˔ ��������C�A������ ��������C�A�����ĵ�� �&�������C�A��������ɚ�D��D������� b���n�u�(��|u |)�����  �ခ���4��� �� ƔJ���%%k���������������}�*���|�*���{�*���z�*���y�*���x�*���w�*���!�i���� ƀ�P N� 4n -�K ���e;SWn �� E�pJus �խHt�c�%\�� �AP�CrR� 0             	 ;HAH�OW�_g�n
� �	�.�/�i���.�n/�i���/.f����.�/�i���v.&u/&����u�.vb/�i���l��� �	�!�������w�!�i�����x!&�����y�!�i���͚z!&�����{�!�i���ۚ|!&�����}�!�i���ֳ��@��b���� / 3(,$���� $ A�<8w3/w+8y���!"f����"�������w!&"�i���"�/����x�!"f����"�������y!&"�i���"�/����z�!"f����"�������{!&"�i���"�/���|�!"f�̚�"�����ך}!&"�i���"�/������v'�+� D. b ��l�Ub���3x�,x�$x�x�xsxcxU s  H �t0&���0�Jt0&���0�J&�/�'��(�'DbȀ�6 ��c�@�� s1!b~�&�.�&&t 1� �~�&��� s1!b~�&�/�&&t 1� �~�&���5&����9�/�8�I�� & 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� 7 � 	�!�~�&��&�r�0sb1f�!�. /�ט &��ט.� ��� �&�y�!�. /�&� 1�0�� �~�&�& �����r0&s1&�h!/� ��� �&�y��/ /�ט &��ט!/� ��& N1�J0�J� �&&3&&3&&3&&3&&3&�>&�;r���� 	A�� �
��)��&�@���E��3I�sE�s !.3&.�(.&'� �%.b %�3.b ��. .&�{ !/3&/�(/&'� �%/b %�3/b ��/ .&�{ 2 ~"��l�!�~�&��� �,qb-!f���w�!�i��x!&���y�!�i��z!&���{�!�i��|!&���}�!�i��-�K,�/��� �-O��� �i,�K �L 3�,$���  �  !!⠀� ����� ���)i*�F�+�l����������������������������������D�ȍ��c� )p�)���L	��SRS�@S�c��LL��� 􉍯�����4���C�� N���U�3�����8@@���R�p.������ZE NW\jw��w��w��t ��~ob��s������)+B!*� ���!�*�/��Jȩ��!�*(/�ȯ���!+�(��Ȋ����!*�(��ȡ����   ���n�)���m�)���l�)�Ěk�)�Țj�)�̚i�)�Кh�)�Ԛp�)��������䎯��8 ��� �C��R1��� ���3�3�3�3 ���$,�Z3X ���6��C��dg .����g�!��� ��F.f��f e�'� �    ��/�����{���c��b��γ(� �g(d� ��c�*s@/�b��a� ��`�*q /�_�^�ϳ�    ��?����?���� �]�(��%2%+d�%�] ?��� `!��k \��l)�� 0[�   ����� 	��D�Ȁ�c�)������
�\[��bo%&�%��DRȦ��c�      � 	����o@)����� �"O�����&��&�!�J�[�&�#��DR������8�H  P� �    �$�j�� ���/�����#���$�j�#�(�!�.!!.&�/�!�&�n*&M,6��  OU "�������r�y�����$����!�J�[�&�&�(�i2,�3�/Db���� �     �     �  �����������������Z�oi"�Y������0���?�����&���2/�3�������� ����T��T ���O�W��f��f��f� u �U�����U�e �	L  `� � �	L ``� � �	00�w����� `K � �	���p0� �� `K � �	���u����� `K � �	rr�rr�`�� `K ������y ��&��Db����c��DX� K�0= �� �  U= \�p�)� �  D��$�k /����&���D�� 2Oe �U/ � D������c�N %������$�kD�/�����cN���SD	�R1�DÀR�T �$�� ��� ��� ����k ��� �D� ���� ���� ����k �.X�� ���X��k �.Z�� ���Z��k �.@X�
�� ���@�X
.�k +�/ � �W V&� ���WV�k �U T&� ���UT�k �S R&� ���SR�k �Q z&� ���Qz�k �t x&� ���tx�k �(/�ƴF��ƴ��� @�� ����P (����D�DN�����DQ�� �D�/�ջ        ] ��/��K �.��� ����K �.�K �.�K �.�襤K �.���� �������� ������� �������K �.���� �������� �������� ������� �������K �.����K                DȀ��c�H� 8�L� ρ� 8� T��T � DȚ��c���x`�X E`3&�� ��� Dȿ��c��E �D&��%5�C�;�� D����c��8L�TO�8��AN(E# ��F�O�&� ��$�� �D�/���c��8L #�C� �$�k                 D�/�����3 � �"#f~ "�~b!�&��&N!"��l#�<##s�!�#�?�#��"�������G��A��������5����4 + �G̸����� ������c��c��c��c��c��c��c��c��c��c��c��c��k                   �����UZOUN3UUU �Y w��e �P��6��6��6��6��6��6��6��6��6��6��6��6� � ���7��7��7��7��7��7��7��7��7��7��7��7��7��'��'��'��'��'��'��'��'��'��'��'� �               ��b�jY�iY�hYZgYOfYNeY3dY cYbYaY`Y_Y ^YA՗ƴv��f��f�af��U �	���������=:�!��<=���K ����� .��d��J��d� �    �C  �� H B	 �Ȍ��+ ������s� ����Թd��0(��@�
�

�?ԓ�(���@���?)ԾJ   ���� ���&��'�	�́ ֖E�	��0֖E��BP֖E��AP�O�@ �?p����  � ������;��A����b��c(����?�����J��?���?��?=���K��C�����'��"��c��k    �
�}�to�nm�{|� �
�Ǫ�ת� ���w���������/�������v��y��{���������d8�9��� � � ���������̂ ��W�fѻ@� ���UV� T̍�������6�;I��h� �   �?)�?9=�� ��?�>��� ������=:�*8��9�����TRN�!   ���沠���:Ih�<��?��>Θ�6��&>ΘF.���d�� !��/�����/�����/�������?=��=��k   �`O 3� @֖E� HP���� �� �TV�U��ހ
 F����&�� �?)�.�撆J� �   ���?�� ���?)��J��   �|�A�|�����8��9 ���I� �8���9I�?���b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f=:��=�Aқ  RQ��D֮G��Ł ֮G�� �UV�T���� � �� ��� �����A�����Ӏh��������=�:?�:G��<):J��<):M��<):P��<)=��7 �Ƚ�A���7� ������y������C  ��LD!  ��N C�� �Q�> ��������� ������&�&�	&�
&�&�� ��ב�?	�<Q�
��N���`1�� (
 ��D�ȓ��c��3��DS�� EN(��I��� >��s �� �D�/���c�ǁ4`N2L�C �L � ������&�&�	&�Á	� .���� �&�X�S %�D�΃T�# ��T5���8A	�	8�R2C � ��A3�8N`!�R1�� �DM�P��H0�����= 3^�D�Ȝ��c��3��`e`�DS��NB E��������� >��s �� �D�/���cŔ �T���� DPS�Iϔ C	זD�/���cŔ �T����@�8��&H΃ CYؖ� � ���R�� 8�(�� ��TO�#� DT � � 0�� �   �P����= 3^�D�Ȝ��c��3��`�1� EDS��TC�� 1DS������c��i��&� >��s ��!.��/����@�� �   �����������݁�#�D�����c��3T�`N����T����DL�C	� 0�����c��i��&����7�!.��/����@�� �   �E��D=X�W%� 3^�D�Ȫ��c��3T�`N����8	(�T5���D �	cŔ �T��DS��ϐ� 0C���h����:   ��켔l~�&���   �~"��l�_�_��_�_�K_�_�˃�K�˃�K�K�K�˃�K�K�K�˃�K_������O������O�. �0� 2�zq
 � ���i�������'��'��'��'��'��'�� ��'�� ��'�� ��'�� ��'�� ��'�� ��'��7��7��7��7��7��7��7��7� ��Δ��Šn��,��ˊZʚ�*ݒ�2��r�r��?�@ � 8 
P���v�OSF=3$3 94RWB[� ն �� ������ �� � ; � ���@����i��&� � ���/�7���Ț�/��� ��/����&��&��J��J��­�l��ɜ��     ��/� �� ����
�(ѳ��/��"� ���&� �&��������b���� �b�����"����&��"����&� ��"�k0 �8�? ����@�� �쁚�                                                                                                                                                                                                