����        8 > '
=95/	#	+	' < 6��������������������������������������������������������������������������������                                                                                                                                                                                                                                                       �+&@ٔ�MA�� ���L �            ���������������������(�������^ E �.o 5&5 �@� ���Ѝ � N�6�����?�@@�e�U��j�U� �����Vw���+� �  a 8 ��gJDYNDFAD=9D5/Dck"g "����-,����  �-,���-,��n� -�,��m -,�����煀�� ?-��� ?-,���砅� -�,����~� �-,����-�,����� -�,��� �l -,���� k� -�,����~��} ��-���-,������w� � �� -���� -�,����~��} ��-���-,�. �(?�r�� ������� n� -�� �m -,���ݚ�ݙ�� H�-,���ݚ�ݙ�ݚ�ݎ �@-���ݙ�� H�-,�� �j -,���� 
�-�,��� �
�-,�i�-��� 
�-�,h���� k�(-�,g���� k�(-�,}���� k�(-�,����� �n!.n�/��-,���� �m!.m�/��-,�. ���ݑ-�,���f�ebdb�n��}�-�,�����i �����"����������⦃�i�-�-�,��i�-�-�,�����-,������i������J,��f�������J,�����i�����,��i� ��. ������}㠿��� /��@� �P? ?`��؇N9"(g$�����c&b&h�- �-ɀ,遠���w���h�- ��-,���ݠ��hҍ ގ ޒ-�,.����~�r��ޔ�!. /�����a���������ތa�b!� ���������`�'����_r��}���!. /���΀����〮���瀮����!�=��!�z�<"e�A��?�g�,������^r�����ݔ�]�(�����\�(������[b������Zb���� ��/����r���� ��}���,�����-,���ݠ���`�'����_r�v��݀Y�!���-),������n�`r��y���_�'��݀X�!���-),.�(?���A�o �4i)3�&����?�u4 U �O���W��n�`r��y���_�'�m���V!.�/��-,���݀U��n�`r��y����_r�v��݀T�!⨴�-),��
�����������Yr���SR��� /-��bX���-�n�/��-,����-,��c�Qb�i �-,�.���� 	A�� �
��)��&�@���E��3��S�������Pr�Ob��m����S�R��b!�⨗��&���N�&��J� � ,	�i�����݄����M�f�ϊ ����l ���L/K&`�'���
.���㙍D.��ف�ݰ��J���,������ݚ��R����֙���֚������������������� �J
�
 ��O� A�_����ݚ�݀ �灎��ٙ�ݚ����J�&@�l�P⡚J��J���   ��X���I"��c�b�����ٚ�ݯ����ٵ����ٹ����ٽ����ހ������ƚ��݇ʊ ����w�H�G�& �τ�F�ٚ���}�����&� ��Ɂ�݉E��n�Dr��{v�K����?�����3��3 ��&�6�
.

����   �(��@����*� /������ ����*�&,!�ʀ��?�������  � �6� ���J�C0�cm��B0�cA��J.��
���&��H�'�.����&��H�'@�&��K      0����5��  6�U��AP^� �����썓D��D3����� 	U
�Yc0�0 ���U� �00� �g���������%U&�Yc0�0 ���45U��89U� �� 00� �00� �g�������A�JKU�c�00� �	YZ�Y]^�Y �� 0�0�`00 ��g����] ?��� `!��k \��l)�� 0[�   ���"D ���m��ԃ����݀ ���&��ݘ�J��ݚ����� ��b�m��ٙԢ����?�/����-����-,����!_bU`�!�S�/R!��~!!&��!bq*⠽�_!&*&$^)$t!�JQ7U�rP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!!.;�3