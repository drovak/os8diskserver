����C� �C1 '  	 	 %  		 	 %     :  �B f ���������                                                                                                                                                                                                                                                                 �������7�&��)��/������bb�������� ����)����J�?����*�?����r��s ����0�����0������&� ?�����c(�����&� �����������b�����)�� ��F��p>�w�FGÀ� �@� ����mP���������T����p�2c����� 0�
���`�����/����l�?����*� �!.b�" n	&�
�
	7�J����F��&�B&�(/�?����r�~&�C����!㨸�!.b��s�&�2c!���&��k   ����;���ȧ �_U������� �����l�6�6�6C!�.c�������f/��"�b�&"��b�b���(���(/���!���,����/���餀��颠����0����< ���&��!���d�J���&�/����k�"H��� �          �	�������p%O� ��?������o �i��S���,�� ���r n&�	&�&�É�4	t�����/�����s��s��s��/����v��0�(?�����)�(�����?!.�?��C�����)�>������8����� ���Y���� �� �1Yw��� ��h�H Y�@������������_���������F����� D��!.��b���F.���&�(?�����c����9�)� ���7���q.��/����&��6@./o!NJ.

���&����� �   �ǲ�&�����i���\ �   �ײ�&�/������� ���� �HYW��Wx>�whB1��X�������� � �)
  ��� ����&�"b�� �
��+D�.c���� 


��(���(/���(���H/��"�����"��k@  ��b&!̿����"�����* ��������� ���8 ����ߠ����� ����ߴ��!����;`���X��H���>�w
s@P��� �?������c�&��D��4�JN
��	&	
&�/�&
	7�J� ���b��&��/�����|��'��'��'��'�� ��ⷷv� � �� ����ר/��/�٦�~���X��
��������)��?ꃼ� �    �����������k��@��� PD���_tȢ��p �p�������� � ��( ��,!�������)��"������� ���(�����(�� �瓓K ���|��6��'��6��'��6��'��6��'��� ���|��'��'��'��'���       ���'��7��R�c��ɉ��(���&��)�B�����K��)�F�P�F%���o_���j�9�������X������ @�ހ  ��&��)��) ���"�����)�J� � �	�����������{�	��*�����/��"b��

d
(?��
1�����)
�9�������t����������+�R���)�j�   ��֣ � � ��  �/���������/F�D�T��H�_�@ ���Pt� ��f� ��>�����0�����S����0�����) ��������"������������y���F���� �          �	��0�����������Ø� ��(?��c������9��`>�?�/������v�	��8L@!W�x���k�_���Z"x@1�Ywh�`��'��P�@ _����� ���c(������ ������+�����b���!�⠺��2�&�	&�&	7D�������7��� �� ��l)��  0��� ������ � ��@?ڀ��"�b!�@��d�É���Dܯ�����J��� ���'�� 	  �	i j ȇhY����0�1����������� ������0��&��<��¢��t��D�����c��ǉ�Á�ǉ�ļ�D��J�
>���ھ�����'��ɿ�"�����'��'��� ��  ���� ��� ��(�J�����F���� `� >��b�8p� ?��"�����'��J������ ��Xp@� >b����b֟8� D]#GL?@�]#GL*@��SF`SR��]@A1	�d� @]��8A	�	8�T5R�C�@I]��8A	�8TT 	Q��@�e6 ]��C��	�ST� E	���e `��3��C ˴P	$�@;]��8�N2 E��S�$N�! ]��C���5TXVCm�P	$�@;]�T	�H�8�F;L`!ԕD�RD	�T5@����1�4�8(�z3 � D	�T5R�C�@I�D T� E	���e `LTSR���D�`6�	8�T5V�C`!�� @L�N ��N`UP28VC`5� @݉4Ɂ 	1��@�`6SAR�% ]�3�8X �5TX�M5z c�VG��