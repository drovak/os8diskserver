����  H� �)/. .5-"%2  / ),% &/2 54054  t     9
8
8


22* 2.    <       2'!4   8 v #���������                                                                                                                                                                                                                                $6�Ke�����ř���2�M`�my�����۪��!:�Hg�~���ٻ �.V�h���� �� �� � �� �� �� �   ��� �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �� � �� �� �  � �� �� �� � �� �� �� �� � �� �� �� ��  � �� �� �� �� �� �� �� �� �� �� �� ��  � �� �� � �� �� �� �� �� �� �� �  �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �� � �� � �� �� �� ��  � �� �� �� � �� �� �� �� �� ��  � �� �� �� � �� �� �� �� �� ��  � �� �� �� �� � �� �� �� �� �� �� �� �� �� �� �  ѭ �� �� �� �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� � �� �� �  �� �� �� �� �� ��  � �� �� �� �� ��  � �� � �� �� �  �� �� �� �� �� �� �� �� �� �� �� �� � �� �� �� �� ��  � �� �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �� � �� �� �� ��  � �� �� �� �� �� �� �� �� � �� �� �� ��  � � �� �� �� �� �� �� �� � �  �� �� �� �� �� �� �� �� �� ��  � � �� �� �� �� �� �� �� � �� �� �  �� �� �� �� �� �� �  �� �� �� �� �� � �� �� �� �� �� �� �� �� ��  � �� �� �� � �� �� �� �� �� � �  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� � � �� � נ �� � �� �� � �� �� �� ��    �� �� �� �� �� � �� �� �� �� �� �� �� �� ��  � �� �� �� �� �� � �� �� �� �� � �� �� �� � �� �� �� �  �� �� �� � �� �� �� �� �  ���� �� � �  ٠ �� �� �� � �� �� �� �  �� ̮ �� �� �� �� �� �� �� � �� �� �� �� �� �� �� � �� �  �� �� �� �� � �� �� �� �  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� � � �� � �� �� �� �� �� �� �� �� �� �� ��  � � �� �� �� �� �� �� �� �        y"�D      P�  "                              ��Jtή"Aa                  ή"Bqך"               ���0J
��❚b��b��l��<��t��D������   ��  @ �� �                    �Q
�%                        �J� 
� <F                        �<1��
                  � T	ή"J[                                                                                                                                                                                                                        @ٔ�MAL	 h��vJ                           ` �       &  	  
L	l �                      Q	    ICQ>X�[Sq5ՀT� V�+�1��? U s5;V��G�Y�x',�U�Qm��_ @ ���8o� ���� ?�*�	��[�S��"&"�"�L��Z)A6`@�I��ffIv���~/�Q�PiM�������Q)�}������+&�0��بS��^c�b��&��6@I� V	��ȷ�f�L��N��;�fO�QL�σ�Hc�|�
��!�N��؋�)�(b\�`�LrQ�0�/�@�)�"���*Q)�:� �1D6�%P�`Z F��(D.��l��(��BF�(�K D��l�{0��F�{0J
�
.
�� �{��z0ë'� �����?����yx +� ��L!�����HiÒb� ��"�""c� �""t"�"�L�� ��n�G)��: @@p��n��&H��ؒ6�G9��t��J�G)� �DVi�(/������!��D&,������ii�_�1�_$�W$��J�_��8��!B�$!.%�/���$�J�B&�$�$o���� �H.�+O1_���aB�BI)�B�(�JP�%'&'�"�L�%&&'%&�&�!$⨊� &�& n''&&z0�'c{�'�z�B�$&B(/J@�$/�W�&$b'�l%!.&�/�&�z�'{0�''&'D�'�%�j L	Lϓ`X�N� �_8�L!��Xi�&w�&]��M������JL��v�/$r��j�&h?�!��$�z����$�B�%b $⠞�$f������ �����&�$&���C�*�O����$z0d� ����n�����Y��/���!$�4�b$Ii��VI)��u�d��u����h!.%�/������t)� �    ���8s"@n�Jޏ&�F.�D.�&�/1��n�.����&ď&����K��"�i)��KŒΏ"f�$�����"�r"��&�&�&�fJΰ� ���� �!���.��$ʗ� ��a) �
�O�@��q�"22c�Jk   33"#3!2 �� .JkLO"NS cM���/L��Jk�h���	�   �j)�j)�j)�����{�w�@��vM)*���耀����������K��*���"��iA�����٦�"�N���`��� �S �3�&3)b(�n33&�(�H��Tْ����(⼀�~Q)I���3&  �}�&�� �� P�n��4cH��q����#��cH����n����$�c�|� �������D�d�b��D&D�/O���/�_�8L�!��I��D�/���.�R%�I���JJ � ;a ☠� :"T��.R)�I�\�b��h ���!.a�V��L��É�y0� ��D�J�C�*ZϘ`���3b� �O�$�fI��$&$&@nW)`� ����b�b�j�/Lh��CgC�&&]iu ����\�R���Ji$�'o���'`.%�/�'�z�@���/LR�!L�%�L�%$f� a%���=�J@
�@/@zn

���&7 �� ������
�&����b=�n� n��J����c{{0J
�J.
� >y �(/���(���(/�.��3�%{03%'3�,%}B������JkLi �8_e �����) M	*;b�w@����j)�pBj)� ���jqr"�0b���or� `�j)��K��p�� �v ����j)�Bn�
j)� �H��3[i�<�('&�<�a3���(��)(&(�"�L�)&&()&(&B!'��� &�&�n((&&T)\њ'(&)!.'�/�'�T\�'�J()&�<�3<'#^)[��0 �X �!]i���o^ (9!.�(f�<&��<((<d<�D���   �;�a ☥� :"TF�F  Q�F $��(��".�L�H �H�H�H^�� �##b[(�:�n<;� � ��c9�9d)L9�mH/*0"9[i�h��)gh��� `��4��c��c(����i�� ղ���D$����D���-&J �OM�k��Kh���o��	c���Úhi��f��/  �!����cՖ�M)R��h鄅f ���J�,b�Y�4!b:(& a.!3&34" ��!�Iݑ�(�TՖ�(�3�Ju ��$�{�$�|$�KZ��<� 3�O���<�I��� ���V�y(�M��̛y� y ՁnI���� m@��p�+(T)Q(�3�JJ �-j)�j9���;�?N�A`)�Z)`��w�Z�@��Z_�<<C<�~<�&�㦦s��<�; +Q0�Q�� h	�Kgh��\t1��L�O1�f��J ��Ji���I鍼* �����`)�Tě $z�M.���?B�J$$@�J�I6�%�+���mjfjjfjmfmjfh���hi� gh��0hy�Eg fuT�*����	 ! "# $  Ϙo�X���&��& f�n��f]ÚM���d	L�r�/��H��b)|�F����7�J� B����fl�*(/� ��X� "ԍj.: ���i��6��N��&�k�  Պlk�    �
��b �/�բ�k�    �
օ+� �Ϩ/�L�RIi�Ly hPH�� �4�#�� �y3�G:��M9�L�@(wBR W�I@���2'�l'�<����"(���'&�&���k�   �'�n8�n��6�c5�g��7 �'�'�'�'�R&��'��;<�i�7�=����7�@6<�Ku���f.} ���bz�.o ���m &#6#\� .W �b�i��k3�G�g��w��w��w�g�uo��o��e5�,k�� pL�R�lk	�u �b@�s@/}@/�@/��/��K F�{ ??7?�K 43�c!@�4/�4�3�J�3⤤K  � �k�$ښ��(���>�K�֊�6i �� �
�
"��b��b?�b>�j�L�RLi��t� � �   �!.�{ !X���bDF��P.�0/�!��!.��K      ��o�      ��c�$bbqI��$&$&A.I��$!.'&$&$!.&&'&� &��&ŉ��<y�(,��`/�(����(��Pq�(������&瀂�����J��"��b a,� 4�>4������� .*��F.��,�" ���E�D�� ba���0�������n w" �k,�) ��� >D@ � 8��?�ѹ����vV� 8 �!p@�((@@  �^��A@Si�R��?Qz��F�8#(�V��R��� @� � �(��""P-�?�?���^����e�?$�^��?�/�!�b>�?�(� ?�o?�o�?$����?f�Q�� ?��~��3�<�ci� � F` � >D�1                                                �J&'eIJ ��&�k ��k   �JO��k ��I��%6�J.R)I�V��� ��%¨ �Z��m��BC FG KR WX Z�L�J��<�<'<B<J{  �@ ��#d
 �� �� ��  +c, 0      �  ? *  Z	�K)#   "!.9b^J� �!�%/L!�%�+}~ � �Ob�� �                                                                                                          & �JQ)JP�Q���@H�P��$r�S	;��)�;!_�er	PrrU��"�	 		 �z���		 	w		 �	 r�SO�R	�w&��"��"-�b��"��"��"��"��"��"��#*pf'�bn T_�a����%\�e����lR%�6�P�Z9		 �4^	`s	`�k               z�(�|(�K ���Áz�����
.��bj ��C�t���kr�&|�k'��'�a�� �������� ׁ��.�ೢ&��� ���'8� ��ՠ/�����t������EEb�����)�hʁ����)�oʁ���(��<k�����ҋځ�� �H
��Á\���J��'�ڿ��(?�D�D7昤g�_���e0������P%����r�6+27Q9R�9SK0~����N�vB 
 vw$ A��Uā�����ߧ�2ԀK�q�$��@� @�eYweW �B�~+  �E�/�{�偌�l��2偌����B剌��^�R剌����؊���� `��� ��!�
��{{�(�́���'� �� �3�c��d�6��C��d�6�O?�|3�J其��[��_   "# $ �fY� Ui!��b:(&(T)!3�]��3�/�(��3�-�/�g�u � ��fi�ciMږ&�
O��O��YY�Io����jCG NL ET SF UR <> cM��`�O����٩J���H���٢���� � ! >< "^ @ 	 E FI NO S_ QU XG M% RW BG ���a 0       Vշf��f>us��f��f��f˳f��f��f��f��f��fU>�g��Pdy������������d����Lc�M��c@L��i��J����U'��NKgu�O����&N��L��/�K������J�u�(/L�� �K���K� �/����(��!� &Jk                        vwf !  # $�&C ���D.��&��?�|�Q�

�
����9��C

�
�������E�����Q)�Q)�"�l��6�<(��H��j��y�QS��?��� �FM)+MHF����jF�w��F�j��� ��j)p�+F�"��bjۓ

�
����9��+ ������jޢ ;��zY )w�W n v| vj)���v���B����e���c�4Ժ&��E��v��Έ��hr�������	M���� L T5�Q�4�E3@�4 R0�F��4@� @$ MD�T5@�3 NR �A��A �3@Eb�Q��@�@�S@�D �# �C��@!@�c��E�F2�C@�  >��@�#�2�5����f$����f�Ь ! "  $�M��BL	CF GK XI	��kR!.L�/Jt�!.%�/�>� y� >��3&�R)3�J5�"��l6�'�8������6�5�k�� p��������6��'**0Ɂl6��  0�����f �v�LbRJk���ύ����ډ����ԍ����Љ���ύ����ډ�����č����Ơ�ċ�0��wG���;�I��X����&��&]��k�(� ��OL����|��K�����/��������n�k�1 �
��'��&�k�  I���à  0��I� 7�
���Ʌ R��3 �DC��0O�#�D�V�C@!�΃DPC%�H�U�$��;-���-�̀F� DT  �� �� @�  � �_��1Gyـ� ! "#  �M��L	�M9�`�d����r��&��6�J���;DH OS TU yz�{|�}~� ���f��f� ` ������N�����v . � ��Cj	Q����jQ�����Q �� �   �(?�Ҷ��C��d��6ӨC��ӣ��t��J��C��zZY�! . `)! &fi]��\��gu� �I��� ���4�b���2�"���!.oq�"�枮2b��d��6a) �(����)X��4&��J�"���      LI2�&������O��q�"2�hm�2dS�J�ˀ��J[ I	��($z0��� ��I��!J�$��$�z��@.0/JI���* $q%�J����ttwttw��f ��`���hß�00��                                                                                                                                                                                                