����  �  8  ?>  ?**    ?/? ?=?      ??8!26&766.71)1%1!556 54*464<408-5	5)4#444 2 88 57194.����������������������������������������������������������������������                                                                                                                                                                                                 
 @ٔ�MA � ���L ������������                               �
8@��	���@��p����� �����/�  z 8  ��@ ��z   ���� ����� U�@�!����ߙݮ��ie�a_�E��A*�6<�0-�Ii�#� ݀� w�AA΃~���**bb�&a�+�/�`�-�o_ +f^ &v)x{�z�� q�{z�� y{�z�� u��{z���^ &�n�p)vx�{z�� 
 &q) x�{z�� box�{z��p)x{�z̐��n�rx�{z��n)x{�zܐ��n�H�� �  .p �pu�x{�z㐁��n�H��]]"  b p� p)ux�{z���p) &p)ux�{z��p) &p)nu�x{�z�� �p)�n�u��{z�"��n�&H.���r&�\ |[�l����Zl)&&bx{�z,�B��n�b\ r)|[�l����Zl)&&bx{�zG�B��n�H�� �  .r �rt�x{�z_�B��n�H��]]"  b r� r)tx�{z�qB &r)tx�{z��B &r)r)nt�x{�z��B� br��nt�x{�z��B��n�H��Y� nbp� r)mw�{z���n�H.�]�]Y  nbp� r)mw�{z��F.�Y �.p �rm�w{�zґ�F�Y� nbp� r)X nm�w{�z���n�H��]]"Y �.p �r�v�q �k�o�pm�w{�z����n �r)Wp)r)tx�{z�B( &r)V p�o�q �vk��n�tx�{z�*B( &p)r)o)q) v�k��nu�x{�z@��֎n֞n �p)ux�{z�U�(�n�U   blx�{z�b(�n�T   blx�{z�n(���f���"�n� &p)&|S�l����lZ�lx�{z���(�n�Z &p)&|S�l����nZ�lx�{z��(�n�H.���  bR&}�DQ�Pl)�Jmw�{z��,�n�O & R b}i��Q�Pl)�Jmw�{z��,�n�] & R b}i��$Q�Pl)�Jmw�{z��,�n� &R �nb}i �Q�Pl)��昊��Jmw�{z��,�n� f��&}��QP"l��.�o���r�mw�{z�<�n�H.���  bsk�x{�z4���n�H��]]"  bsk�x{�zC���n�  bsk�x{�zS���n� bsk�x{�z_�움9A�� �
��)��&�@���E��� 0�H>�n�&&s)��d�� bkix��� � �{�z����n� b bs���r�o�Np	q) v��n�&�Z�lx�����J{z��9�nn� bsk�x����D(��{z��9�nn�  � s)kx����D.(�{izד�  @��d�� �v �J
�
��(��H����n�^ &v)x���^�M &}P�l��vx����^ &nv�x{�z � ��n^� bvx����&}L�l����vx����Ll)�^�M &v)x{�z� ��n}�Pl)�q��q��n�q{�z?��nS�p}�Pl)y��{z�O@�n�}P�ly����Sp)y���P�ly��{�z\���B/l��c���� �>="khw�n�^M" }iPl)��vx����p^� bvx�{z�� J�n��n�^ &vx�����^� �nnv�x{�z�� ��nr�^Q" bvx�{z�� J�n�Sp)ry��S�py�{z��@�n�rq��q��{�zȔ�nr�qۚnq�{z��@� �S�/��_b$���������J � ���y�xH.w�,  ��<�Tl�Q_f�n�_�&Sp)ry�����qi�{�z ��n_��Sbp}�Pl)y����&q��{z�P�n�q���֮nq��}�q���֮nq�{z�$P�n�^ &vx����}֞^ &�n�vx����K n֞^L" bvx�{z�8 Z�n�^ &vx����}֞^ &�n�vx�����^�JM" Pbl�vx�{z�X Z����W� �a�0�n�^ &vx����}֞^ &�n�vx�����L�^ &o�vx�{z�� Z�n�}֞n֞L^" piv)x{�z�� ��n}��L�^ &�n�rv�x{�z�� ��nq����}֞no�q͚q͚{z��P�n�}֞n֞^J"M &Pl)v)x���n�^ &v)x{�zЕ ��nS�p}��n�y���n�y��ny��{�z��n}��n�Pl)�^�MJ" kiv)o)q) r�v)x���n�^ &vx�{z�� Z���n�^ &��b}i&Ll)�Jkv�x�����L�l��v�x���خ^ &Ll)vx�{z�" jπ��ƄI�b�&��
I�b�& � ���J�� �+��Z,)�+�[b,��+��\,)�+�]b,����@	�0T`��&�n�&&}L�l��k��J�n�^ &&&}�Lbl��k�vx�����J�^� Lbl��v�x�����{�z�� ��T`�T@S P	�T�@��C ��T` �	CBLT@&XR�� S�"��3��@��T�` M Ք3��X�D1׋M��h6-���C��ă  ���n�&&}�Lbl��k�q�����L�l��q��{�z ���nn�bSbp}�&Ll)�Jky�����JLl)�Jy��{z�p�n�}*�Jp)H.���  b �noo�Hl)kx���� x){z�@�x�n�}�H��]]"  b *bGp)�o�oH�lk�x��� �x{�z\����n}�H.���  b`ro��o*�Jp)Hl)kx����`x9{z�y�x�n�}�H��]]"  b`*rGp)o)�o�Hl)kx����`x9{z���x�n�}�  b oi*J"pH�lk�x��� �x{�z�����.��$�&�Ѭ�qYNa㳰�N��T9?BQ箠S�jl�;y�$6��uO�g��=��8n���/��r��ޜ�. Z�� (�n�}�  b`�~o*�Gp)Hl)kx����`x9{z� ���n�}�  bKr *bJp)�o�Hl)kx�����n�}'�*G"p� Hblk�x{�z����n� b`�~o}�G*"p�Hbl���� &kx����'b kix{�z=����� �                                             �n���[&[o)}r�6H.���  b*rJp)Hl)��r'kix��o)��F�/���{�z�����b�nn�}i*J"po�  fHl)kx�����J�n���b  �  &}o�G*"pH�lk�x�����|�Ob oiHl)kx�����J�J{z�����n�*p)H.���  bsH�l��' b((bx{�z��nP�*p)H.��� �no �sH�l��`(6(x){z����n�*p)H.�]�] & s)oH�l�� (& x){z����n�*p)�o�H.�]�] & s)Hl)�`�((bx{�z6����n}�&&*J"po� &Hl)�� ���b kix��� � ��{�zO��􋀟�LV2m�ح���:���n�*p)'b  bsH�l�� (&(x){z�����n� & s)  . oi*W"pH�l�� (&(x){z�����n� & s)  . oi*P"Wp)Hl)� �((bx{�z���Ƌ ��n؞*p) ji�n�}H�lh��{�zǙ���n}��*�p ��j�Hl)Hl)h��{z�����/��#{8���	�����|�|�T���_��n� & s)  . oi*J"Wp)Hl)� �((bx{�z ����n�  bs �  �o*�JP"Wp)Hl)� �((bx{�z����n�bbs��&�J &&*p)oH�l�� (&(x)���� � d�{�z3����+�/�޻���n}��j�] &] &O&G*"po�Hl)vk�x{�z_�������2;��� ��n�}b��+bEc�bH�� �o��!�⨢� /��I Jp)Hl)kx�����O���D�&�{�z����� � &j)�n�h��{z����b bji�h��{z����a��gҞcg�^���f9g`� f)gr�,f)�66�O�g�d#�f����gh�%f)gl�'f)gf�$f)O�&�����ZCր�^ ��n�}b��+bEc�bH��]]" oi�!.��/� �����IJpH�lk�x��������D"��j{z� ���n�}b��+bEc�bH�� �o��!.ƨ/� �`���IJpH�lk�x��������D"ļj{z�.��݀��n�}��j]� ]b Gb*p)oH�l�� Hblv�kx�{z�^�������!?� ��n�}b��+bEc�bH��]]" �no��!�⨤� /`�I Jp)Hl)kx�����O���D�&�{�z�����n}�b�&+&E�6 &�!.¨/� �  �IJp�oH�lk�x��� � ����D"��j{z�����a�-`'cg�ۄ�����nꛮZ�͹W�:�\x��+9�����w����v�z  fj)x{�z���n�  bj��hx�{z�	���n�}؞p� �^ &j)Hl)hv�! ⠭�,x){z����n�}؞p �ji�Hl)h��{z�6�����n}�&Ll)�J���L�l�����n�}�Lbl����n����� ���� ���� ���,�,�+� 5�N ��`1��	��9 ���6�����������d⛀cIc��CL����R0B�& �g �cg�^��f)�D>���gi`�����e) f)����D.���gib!�e"�f����b��bAb�b@��D����$��Fg�f9��J-`'@�⳺D����D�J d"   t����DM�P��HG1L*�����ʇ� �C�&�ą����q�� �))b! ⠍� ���R!!�/�"�! ⠕�� ���#�#�+ ''�-�� &&�-�� %%�-�� ���� ���� ���� �|�Pb[l)�J��Pbl����Zl)&&b� ��l�Zl)$$b((b� �|�Sbl����Zl)%%b� ��l����� D |	&Pl)�J�Z�l"�|�Pbl����Zl)R!� �b
�_?d�_?d�� �>d)=d)d�� ��<�&�_ ?d)�.�晴J;d)� ������F�C0(��@�
�

�d���(�:�@9�;d)��N���� �&!��"���� �S��v�k���&[l)��J�Z�l&�mu�c8���KO?0 �l�l��� ��[��-`'��6��������`.�k��D� �   E�67�,65rQ4r3� ���n�b�}i�� �Q�Ll)���D�懴J���ԟ֭&ՠ&��6��0��'��D������W=�B3�-$�9F��NĀҀԀN�̀�D��C�À^�T@SXGS�TR���@MN0 ���R��C 	�H��HGS�TR��AX�K@��� 0�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C C G�S%�RA��DτTՃ�8��C ��NS��S!�D�H�4Tn ���7��� ����    {�����