����@  B H� �'29 1>+$'+''+/  2/<'/  >   ? }1?8>* 
?? ?&>*7>222  ���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���������(����	 ���i��@�
 �
����'�'�&������#����P����	�bc	s	s�	'	7�J��0��s����s��s�n .��s�i��7�a� ��y�nƉ������y���H������ TU�����jh�������q���������w�� `� ����2!@�/�����!.�/��F���&���K�L����Ɉ ��
�"�n&�����&�����c���Á��ӣJ�����r�j}k�ެ�������ײ����r��{�5�����+�� �  � ����
�c�
c
c�
c	
c�o?	�t㉬
 ��?����KqI�����/� ��T��j� �����������������m-����ˁ� n�����������r�|������� z�������s�/��F��&��0��&�� ����� ���|�"( ��/��¨/��"�k娟���j¨/��*瀀����V��8��������W,U,�@TP#�K�G�ۧ � �f�)
   ��(����b�b������c(��F��2�l'"���O��rF�''�"(��n�|������ ���b�(/����"�b�� ���(�� �&F.���b�Β�z � F�����k  `   m���U,d�lu� �S������  ���?����q>(��(������c�(�F��N@����/��"��c(��� ��V.��c��F��?�����)    �
������r(�!��&��������'���L�O��"ʁj����%�� ���j������bF��"�c��ǣ�N!.��z�O��T��p� v�������4� ��������'��������X�����������������'������� ��,��y�́̀�遦ʁ���� �	��ωp���������U����
 �	�pĉ�����ư�� �  ����"��c������!>���� �À���:����f�m�o��j�T�[A� ������ ���cJ�����"��r��&��; ���<�� ������i� ���� �� ����������  � �H/�����$���� ���췁<c

�
�������J��(��(��L� �(���@/��&��!��� �jk�"!�ہ��(?����C�(O��牬��{�	�' 6��JMT�� �n�o?���V��?�������FN���&��,��|��C����������i�����i��������(������H@�&���� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d��������D��� ���޴� ���� �&�&� 6� �bk��� /w���,m�ڀ��	nj���� ��� &�&��K� � o��b����)��i#b��##�� d��H������ђ$�n%�j     � �                                          �Ty\ �T ��/��釠�3b46b75f������3D.D�@��%(/�������5v$�/�خ�5��������r�؞�s����@������Y�$�(��H��)+&()&'(&&'&%&&5h/�����5�/�5��n4/�4����4� ���3� ��퀾�)� �   q \��L��̺���?DV@���]U�= ���  !%f+,&&/&'�&(�&)�&���@,�++&��))&��((&��''&/�&&&%�%�h%�)�J� �$�/�ؾ��5 @������ +D+�).)(b(�'.'&b&�%.%�k �            *%b@H��%&b&�'.'(b(�).)$d *���+�k  ����`�� GE�N,�������� .:$f%&f'(f)�n�:d�����7�4P.(��@a�4n���n� �4�J���ܤ45&��H���ه��8�!5�4�n�Μ������S��O������'��'���� ��4���J�9���~�l�ܨ/4�J   )a.)n(!.(n'!.'n&!.&n%a.%�k ����Y�R  i�� ]�                     S �$�$�i�����߅�.%U//%*�&/-$"$o.#*%&Q/*n&o/#%(�	�%�o���*.*o{��$$&*�/{%�@���$ N�O}(�$%fQ&��/$(/? ��?�   ���.�Q@��}��O%.�%Q@��}�� %�%�      */�)�I�$&��������/�%*��-!.$$&)�$o.}+/��/��*�@���$ N��{��!+�/a.+/�+� *�*�n+(/��/��}�� ����%Q	(�$%fQ&��!�$$&�.�%                                                            ��/�)�� �.Q}.�A/�������.��?�%�/���.Q%�j-/$//H!���b��/ *�Q�Q϶Qo�$b-Ƴ �Q*��%�*� Q �#*�%*� �����%�.�/�خ+)/�ڮ���	%�! �-�$Qo&?k+/�%�j                                            �  �/�͐z�F.��o�<��t�����(�����r��~�� q    !ϥ���?���D����&��!�ʀ���(?萦��É(��Φ����&��&�� ���9  �ͣ��I� �
����"Ͱj ���&��2@������0��'��J� ������� � �x�?���������������                                                                                                                                                                                                  v       �   ���                    �  �� �                                        �                 I� y4     V�������0F	 q�*�=���c  ��+��/.
 A�5? ��a\ �� T �8� ����L������K���������������� ��   � ����  ~ (����!.��/�����޵�ҷ�cH������v� (��� ��B���� �����H�� (���b���)D��H/&����/�5��&�b�l���Jj�����T���7�- Ww&63��9�nӇj ��i��̪�̪̱�����?��CH�(� �����̏�!��"�`&��X��j��},b�H.�����;�/�ӢD�� �����	��}�
�̳����D.Ҥ, �    ���l��&�����rD�₁��˒�'��&��& �&�|���&����d����'� �   �� �~�{ �zіz��6fy��c00b�:f�0�x�����/u�/n�/r�/c�/������ �/� �/�9�:b(� �:dw ���� � ���ɼ �0H.@��n�)�o0.��� �:F.:D.9�*�" ����'w�/�&0':(/!��w�� �����/v���������3"[�(��"��h��u�����0uI��/������� ��/�u�t��s����r��bF��⩕�'�0ē � ��� �:&13f2b���"���x)�����f����� ���������������� 	 q	����p��q���:��!N6�n�j�����:&����gp���)�a�� 9�9��@.o/������@O�9����9�c��o��� n	H.����v����%�b&�h��sV��s��m2�t�y�!.li�Ȩ��8t���� �
�

�r� H.��&��!8���y����H�����J2����L��Ɉ �
��� �� z	w�NziOkiN� � �6d3G$0 Ə ��j�i8�`o�����H/H$.����2 H��2HHb&��8D.8�"
�k� ��H����H�HBbhC�D�Fpk��H$.����H�HFbG�h
7�Jk� ��<�
�b�b�k �t)@�/����t)C~ D.����k 8F�8(/��"<�h
7�JB| �J&@�+�����?��:{ �@�/gھH����C~"Ih!>FF&p �`F�Fo�C�f����$����8��eb��kU�_CC4 d���/p����Bh !C�H���D��Cf�H�H��H�nf���тDDb�/�C�C�i�Ѩ� �Ch0�CdCh0J
�J.
��                                        � (�p�o�,&�n1�j�2�3�y�4&1�/67&5li���c3rDD��&%(/�ȯc5�$�/�k��n5�*�k��wr�k�s��2�/�5�7a.4/�4�3�n� �7!.5:&3�/57"5cc���5h/�4� ��!1� � �$�n%&f3�/5&5a.4�/2�/7"4@/ ��H$�!��!��k��d�֫    @ ^�h U@����c�X�$�(b� �@a��&�+%b&5bh���1�������5�/�5��n4/�4����4� ���3������ �t:�@H�1:�����:`"H��:d���`"����(:�(�2�(��3�b������֮݀�_)� �+�j^t)+�J� �!�+,&&/&%bib.�]b�%�(�J� �\t)�������� .:$f%&f���sx��%%���.��-��E��"��0� 	4�d����/�9��kilע�4��c�:�JccY��J74"P(��@�a4����&k �4�J����פ45&ccYks��i�8!.54&k��� �        ��1�/�5���/��+ $���k�5 @� �!��t)�J� �*��?��ds���	&�js��n����^t)�s�x����_��_� P���H%�&n$d�y� .li����)%�/��"t��!.b���"H���n���*�j ���s���	&���t�� ��eb�! �����| ����b
hb�o�<
�t�e���	����;�K   GA���V���p �H X (	�H��(��r�^&��@�"�����h
o��n@�/�@�dx	�L��4��.��N��C� 9m@/ԗ��	�w����!.��0����\��	�	�n&��(�Ȗ���|	���	�h�
 ^��h �	tԼ� �� @ޛ �����f�IC�C N��� ID�K�D��C�C�d���ѓ 0� ^@r���&�/�֮A���xO��Po�Uo� `�@���/�o��n�b9�n��&@�/��@��9��������؎Ɂ���CCt��
 �F��Cc~C�h CC7C�@� ��J���&C~ ���FE"�Bbh�Ga.F�/A��@�    ���F��C&� �� p  	� p yT �w #� w��u�p60��{ ���&�@b�g�y���� D�Bh OBb|J�H��N�jkN�OODOyIH.���D�J��/�p� {	 
#jii�8$�F�
(?N�
O6kL�݃* �Bh ~O&�I(OCv��fI��p.O�<����{� j)i8�!�jk��ii88B�JF8b!
�jN��
'O
'G`.F�/�H���~�> < U�z�w ��&z��| H��#bh�#��/��!#�##Ch�#|0�#d#�6##C�b(��h&��"ѥj��bh���&��| ��b!(�hF.4�� .@���&J.

���&��)� �   ��"�b!�� ��kߗ �       ;  �  �  �  ��� v�    P     P P�����z ���
��]��Z\�X(�@��X��  �  �  �  �  � �ko� �Ƛ&��'�8&���gº��f��(ܵ�|t	��(܁���<Ф�	����е���&�%&}�(%�J�J�H&��y��{%�%
.

�r�%r �Ћ ��"�b�t)܀� �=���ky� �� ps �+��@�6#G <@ d�2                                                      �            �             �            �    �                                                                                             �$@.�(/�8���%�*@H��8�J8�k&.�%����'#"&? �+D.+&b&�%.%�k  *%b@H��%&b&�$ N*�J+� �&a.&n%a.%�k @,+"+n/&"&n.%"%�k  �����& ��P�#[boڂ��o#?#�#O���J? ��           �L,�υ�	����[�)�9��	�Y��i��i:�y��yE�i��t�y���� R�SRQ��� 0�D�8�8E ��T��C NT(��C N ER���CR`ob�R1��D�8FN`� 0� R��OA�R��D	�` l.�σG� � 8�R1�� � �i � *jS�F�W� |���+ �FF&D.�f�� �����
&

C  /�
���w=@&A�nqi0tiu0� ��^�+kT�%�'&�'0[b�ui(^�t0�ҵJ^t)e�&�F.���.w�	��Jq�����kk^�     Rڈ \�  �  d* �o�A� ����  � v� X v �      �����A�~                                                           �o�%� �8�k ���Ɓ���J ��آF�Ǵ� `� >��b�8p� ?��"�����'شJ��� �� ���(� � ���ឋ�?� � � �ƀ � (��!��&���Ћ�����������H������� �� ^ �� �Ŧ�   � 5`DR	A�� �8MRQC(�U �!8��C ��MAV�C`!R��OC�H�`1�UDRD! �A3�8NR��� �TD	! P�TO�#`�� ��6�`   �@��OC� Pҏ� � X� 0��� �UP2 � �RE �@MG ? ���� �&��6��� �d��'?�� �b��{   Z$&#�&&bȠ�%+f�/�?�#�&�&�#�#n��cJ� O�����O� ���{�"��n�㶯j&#&%)�k&/z�#?{z�#�:�/���i8�����&�J�����n�ss"��&k�? �v �     v �� ���L̈\�c��z�F.@�w��&/�D�}"�@"/��@�w##T.#""#n��o#�6#O�#��w����&�&z��| (�����&�@.?��D����)�o��* �����o��+   J�!/��b�@P��\�މ���k��bX�Uޕ��q��`������_ݛ������(��ۋ&z#�)�l/� ��ϡ�w@!#&��6J.r���&�!���'#!&?��J ��|J��c�%b ��&�/�?�# &���,��{|����?�������������Հ�$�"�?��۫���  ���w��{HIݟ ��޷�	�֖�?���һ�ɤ���U�\͜@�Y����o�/##�?$�-b�$��w�Z�(#�!�$ .H��a��?�-$&?�Y��J� �#�b�$f� �##c#O�-�#.6#O�#�/�l�����'(f)�n�j���"�rH �F���'?�����+�]?�##c$#d���##c%#d��#&6?#�$#'#�J�#�%#'#O�&�#?{�c���@L�                     p �$�$bi������$�$�f,%b�$��.�/�h,&&�%&%.���+�/&�J%%BH���+��Oc%��$��/$(/? �a?� ��.b����۔/D./.b.�+%b���c۔ -�� � �-/b ��+�k/./o�,�&,&%��.�,b,�+.+-d�ܫ ��H�/)�I�$&��������!$�$.ba.�&�+/b�����&� �%."����,&�%�%�%."%��&�&�,�J�/�,/�@�&.,/b��a�&n,q.%/�%��+�@��@&��%�&.&$d %��%��&��!�%@n.%"��% n++&�%�(&�%�h&a.&o ��               ٵ����/)� /a/�.�a.������.��?�%�/�$�a-�`��!��@����(a-�$]i�?��@/���a�����? � *�.@.H�.�/./-d *��,�k %(&�(+����%� ��&�/���YȚ$+f���%&f� �                                               +,f���/�                                                                                                v ���s�/������r
�b
c�t�����k ���r��c�/��
�b�j��� kj��          �����E� ��fV��������U                                                                                                                                                                                                