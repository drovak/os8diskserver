����   �  �P P  � � �  .    -02? # 	 /8 	 	  	?   ?  #  . #�������������������������������������������������������������                                                                                                                                                                                                                         ��ʒ4                                                                                                                                                                                                                           �o� $                                    g�"1 �g                                                                                ��l�>F!l��(iib�����D������F�!�晵¸D�������F���Ķ�J� N�F�ȱ�$��+),������      �����b�����c��   ֌l��&�� ���� F��,��   ��y��� ��6����s�!��/��� �   ��Dݑ�Xi�ę|� �    � Ã2T      �:0��b��&�{0J��4�'�6Ù����6�� ��l�!>�������F.��)H�������D�廬��4���s
����"��sY��A�����������6�X���r����皙���4�p�l�?2 �c�op�  r� &p{ }����+ �l���   ��no ��@D�P\lUk _`8U2@]EUX5U��b~���Xn � pr��l��2 op '���ÄT� H                                                               ��!                                                                                
 l�                                                                                                                                                                                                  � �������������B B   12   -   <.	2$??????    > ;< "	02$1  .  ?:            ??            '8
<(*5'?('>; 
)'=
&
(
*
+"	
& =	5+0; '
)5-8 .-  '<"	                                                                                                                                                                                                 */';:9'8'7'89+'6.?8        ?-E "*.058
)/E64		"60&! F   	    
    1  " !2   	 !  ?? %       -   	37   ! !09;   2	*		"
"2 			    )    	   2	:		2 
29 2 2    
					/0G;H                                           ?>    /???                                   
 ???  ; ?>>	==><<>;=;:.4  ?;42/  $,9$$  $-$"+> +8+!$-$#++76(   ?!+>(/#'8+$  5?'4; (I1I4-8	# ,+*)(�		,5/   <<<?38;=?!??(?< 
      ???�����������������                                                  ��Ñ�ǉ����r��r��r��r��r��r��r��r��r�|��'��'��'��'��'��'��'��'��'��'��'��'��'�����'��'�����/Ɖ���'��'��'���          �
�K	�L���6�@qH�< T 9S�83�7�g�tf�{eYw��IW�|Z3tX�|VKJfIf~l n�\2q@ȁ���<���������3q�b�����'��'��'��ΰ�l����L��)�,�|�!>��/���q�n��l�7� �4¹�la�#�o�R0(��́��D����<�G� ���F�!���&����J��&� ���K��CT&  �                �� 	0=�<EPS�O3�N��*Ñ2Ā|�-�<-�~ 3� @	�L�O� 0� @�N�� 6� @!I�i�i�,�����<m�bm�&$ړ!���`/�����| � ���U��Ñ|ƃ���c��l�H.{����:���&��'���� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �j<�
�  ci| f`�P�m� �|�,�����<uucH��u�}�H:�Łl��<ddb��&��?������dD.E4�db:5��c��&��ǁl��0���Ǩ/�u��4�����F��x�����      ]��l�,��|�� ������J���{k�rF�=��`"����.Ȁb逕��bC��D.��"���w�y@ݟ1J�}Dp�P�du  ����*��������$9���ˁ�Ñq�q .��n��ni,i`�&�i�����,�$7�i*),�����i�D�i�;i&��J��j    J � -�-Ǡ �7�  X a2'��ĂL� ����l���ٚ������à����K '�g Pe�\��������� �; ���竆�2yr\Frp���5�Dq { ��l�&��BF���/� � �}�ƙ~,��,� �$���!ɮ�����!q�����˰�,��Ƀ�˃�� � ��Y ���=0`�/�Ǯ������|D.�������:0��&��� �� ����k�/۠���b���� �                            ����)�o��`8fEP����	�;����
���� ������8���  � %�7&�(&�
&�	&	
7(�J��2�����(���P.�/����4��%O�(o�)(c)��)�()3(�z4��� �%�"((c(��((b$b	%bH�!)�!>	�?�)��(��ϴ� �          @	Ui% f_�M�T��;F                                                                                                                                                                                                 �<�|�/                  ��"4 " �1�Q"�8#�Q3�m�                �� �� ���s����   ������      ����               y@� �߇X   �                        ���������� � p(���H� � ���¡�f��&���(���/�����J��#�����)��������)��)��������&��6� �   ��@��������&�������¢���l� �   ����&�����i�����É����9��'��9����F.����e������� p��K��� � � � 	!Q67�>?^gW
�; ���(����ˀ���� ��(��(���� ���b��/��������(��"Ȳ���"����� ��K�ǎ��/�����{��8瓋�  v��PH �   ��㾿d�
>

�;�;�� ��(��H���(� �&!��"���� �������  ��(��(犰�? �@��H���{ހ����� �}��  �	��)����˂�  � ������������{� ���c��r����!��)��%���� ��}yo�mn�  ����@O ���6��&�Bl�ͿJ̿J˼J��L� �    	�YBY9Y������ �� l����b�����۔�,�|�� O���� :7�9�8gW
   �8�HT P�Tq	�SN��E  
@��N�Tυ��@` �Mp IC�
ASUN Σi �Mq�`1	GS��%` ĉt��T�C�D� �  ��qVS!ԃ킕 L� �4�R@ XL ##� p�8vV�C`!� ӇLC QV`!�DE5� @�LqC �TR�MTR���s��D S !T  Ň�8�� H�D ԇS �# � H��p�8 ă`�`@�� H �R�  XS� T� @��c] NT" �@�g�=8 	� ` R�$= �S� `_ ��E@ҷA- � �N  T` R�� @τT �  Pσ � ��� ��,.(���� �       ���'��l��� �����6o��������/��������/��������������������P p���!�扮½�c��d��6��B��b��l�?��s�!�Ǩ?��� ���D������>"��j$Г�Q���$Փ�$��q2 ��i`bgid�i����g�J��J,�����iB;�*��C��@�� �q ��"����l6�m6��6�l�B&h6C��lʄ�Q��Ũ�$'l���x����-Y�$'����-��m�*-�-h�����/�()-K�(��+,��j�h�/�Ũ��� � �i*)-ś ����ʻ�C��#� ��8�L5`I�C � ���X��4 ��8 8��o��� ݦS1Iw��0pm lR�H����·�.6sX�<��2b��i����ٍ���r�����Ȅ�$딦+),���  i�Li�,����B2h�cn�co�c�߸��
�s v�!9�F���̘�6�6��3 ^

d����6o̣� F� �� �|� �����c�o����|� �$w� '�s @\�h�y�)��p@on ln�D H����Y0��s
����"��y�A0��~��y�A0��&q .��b����Ӛ�E0pqbD�!p⨮�p>"4p&�?2 �c�op�  r� &pE ��bH
���& �0� 'p�&�X� ��� &p� �r>�&��J��Ā �� �s�� \� �q .if`g&�㸏E X
l ����n�op ��@��U  �    q  ��	&4�&��	�r>�& �J��&��&ߘ���	ǘ>"��d�ߨ>�&�	����>"��b!�⠲�4�&��J��D�q� ���	&��&��!	� ��>"��b!����4�&��J� �����b�@n?��׉�� �q .��b	4b� �                       ��?n�P�� �f�b���ccbG���6 6cE 4�& �̉l�� �(/��������������� ��/��cb��b  ��b�k�� ����= ��&�̲�Y����= ��&�̲EH
����k � ,�?(O�)_� P\�i������Y �K()�E0H
�*-�� �.\�5[� \Å?kF)f�� �a7�`E��  .ŷ�ũ�����������Ū��������������������¸jcD.E�4�&b�bƷc�����cb��b  ��� �  Db�h �O�쐴�c.�b�� Ǹ� �cD.E�4�&�-��-Ǡ �?��<b�4a� ��˒��;;R��&!ܚF��i���;H��6 ��"��{7 @�I� �Q	�t��U D c `�P�`TR�8��0�N2E.X..� ���CC��  �C���$�L@M������ 5A5!�(Ձ��`XN !`DЁ� �8R����@� @���NTR�ES� �S	���D�MAc ��<f�����C���# P ����_��2XD�ԃ̃�5�T@`c  ��e�����D̓ �� �   ������P� �� ��  ����l��&��?���$b�o��'��'� /�����)��)��)��&�.b�������J����g��r�����b�(/����	�;33C`3t�J��U��� n
�i����
b���h����
���|���g�JO`�gib;i&�P�z'��DNKw �      �? �@��� �� ހ�(/���(���(/���(����t�����c���������(����/����֨��(��(�����(��(�����8� ��O�&�B�!��"���� B�������+ �����֋���o��K�����|��'�֨����K��'� ���s���A )w������}� ���"��f��i�O� ���"`��/����D.̯bH�����$����"����b�����+      �r�����/�բ�bb�b��c��������&���
  �β�{�	  �"����"���"������B��AֶM����T�{�<���	�������	�� f�b�n��f���(���/���" ��(����/���暀����"����H.&/���t���������&����"����?���h�����h̀���h�����)���6��6��C麚 �	b�ڛ�����빀��� �=蛮��S����?�	���A�]�� ��/����/��b�c(��(��������︻����6��&��9   �
C٤�@����F����������D� �  !�(?�����D���T���?��?�˻���^����@�(����i�=��ߛ�c�/?�ߛ�%� �   �^�]T  �p���� �N�]�x �&�(���p.oN�� .�{���@�����P.�/��K���
��&�&t����ǈ�(/���(���(/����Ǹ�����(���(������<�����&�����F���|�"(���k ���{���#� �-��pߧ�W� �`��� կ
F� ���6�������/� �� �b

�
���(� ��(�������� �����������(�(� ���i���������/��������/�в��(����/���!��&����̯k ���4�l�<����<��@����/�ԋ    �����ꋀ��!����}] ]��� ? �M� +��������6��)� �����)�������cb�����)�)�)��� �	#�� �	+�� �	3��r:��:P�: �4 �T��G �J F��: �
   � p!����N��NJ p���l�׊��(?�����������ݺ�2 ���J��+      �` �� T*pL�K ��� ��d Z �	�� � ��/����ŀ�  ������ �	� �� ��6��'��)�&� ���4(����� ��b ����É�� .�/��� ���(���(/�����ǉ����  �����i����� �  �������  루��  ������  �	 � �	  ��D�p�������  ��W�ͳ� �	�����涃l� ����H���b��i��/������.����@N��,� �� n��&�����0��d��0J
�
.
�� �    ��C���P�`�V`V�`�Li!�`�`@��k�R� �������ҋ ��|���ỉ��w���+����8����� � ����?��p�T ��'�����  `         ���� ����� ���c�� �� �����e �줈��  �¨������ �$�����+,��� ���ǉ�� �q .��bqbD�
�b
'�B
@/Ҁ���Ɉ���$��������������#�O ��]g0͎���_�O���y�����-�<-�~ ;�� �\ i-�� \�$�����qb ��i`bgidi�,�����i*)-��,�g�J��J��˃i�;�*M`�d��4�Ӄ����C1 ��6�����(��Y�&�:05�&��2��cY���6����'���� ����[� �   �J�
����+�H/ �.���+��l��=���� ��� ��6��N�6��C��d����d�/����<t���� ���˛��E�����<���O����:�� ������7��������&��2������� ��
>����&۠?���
     �̲��r���۴�(����Ͽ���<��~��r��r��r�G������������� kyP�]��T� �(����bF�����b��&��É����)��b��,�ޖ�J.����b���݁l���JP�����P��"��&��"��c���@������"ہlۉ<àn� ����B��� ������)���Z�������@�       6� /��
�  ��߀� K�NjZT�]��f�hg��F���� ���?�������FN���&��,��|��C����������i�����i��������(�����H �&��� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d������ ����� ���� � (����B���ǉ�� ��������9��s������C���z�����ɀ 5���K(����� 5����� ���s!� ���)��)���F�����É ���@Ŋ����f������{����?���d������L�����ѝ      �ʌF��:�?߇( �TN�<0��?  ��/�����b��b��g�'Ӝ'�����y�&�|���xD��r��'��c��������Ө?��0�����0��s(����tĠ?���������������N �	���(�����<H����)��+ ��bg�J������|؞� �-�����N0 ?� 8G ���Џ���k��ߗ��                                                                                                                                                                                                 �;��V�            ��  6�	$��2��"��$ �o���f��f,�t �D �v��f��frdJ'uIG�6�  4N   	    8 ?@ �� �� �� �� �  �J`HP`��������������   � �� �� �            ���   } � � |   ��� ����	�yr�k� ��� ��$������$��!�F���c$�����$ԑ!��F��g�$ݑ!��qnqD.qt&qC t .tqb� ��qr[�/��������'��'��'��'�Κ��'$��Κ���w�$����᪠����{��{ � � ?� � @  UV��s���f�O� NWY��,,�q�/�$��������$�ٌ�����'$�ٔ�����'$�ٜ�����bԠ�����r��r��r �࠸���'��'��'�� �����'��'��'�� �����'��'��"�����'��',�          '�a2b c���K�����������̗6���LT3R83�A?�3�%3�3�� �� �4�l�	6	
6	 6 � �|
�J��Kq�(��!�ţ& &�	& ?  s�!� �?��� �	�JO���>�&�S�� ~ �◾k `��'�)����C��#��V�SO"�c1�A�  ���P��Є���X E30-��@���-?N x������
�s v��8��O��  ^��/�#@�À^��%L��qb �����O���� ��()��  �)�= D�iib��)�����b=���c��b(��D�����Y0l�cA!
ib4�)��J`�&iiB�њ�i�
��V`�
pb���ĕ�� �#�V�����  "  " o"�
&m�)�l�Ub!�l!t�@�W���cM�[�T���B���L�(/������ �             �
���������(/������ �             �
�Ū���Ś�(/΂�Κ� �             �
�ߪ���ߚ�(/났�� �             �
����ރ��䳑���z�������xwf��x���f�ndl��� ��	&	�6�eb!��Ș��!.xf"Ȗ����/f�&'��	 �o 	�	c���	�	d	�6�G���t��������EҠbD�E4ӠbD�����R����d�bf�b�����lH
���;�"
 n��&��
�r

w���x� ����d���         ��rxb(g�h��}�g~bh�j&(�2�?2���B,���� ��������bn�c���(���c��lH
��ƟD.E4�:b�5��c&���rw �����dD.H�E4�db:5��c��&!�Q)��cr rbr�v �t�A�����!�"y��X�a2'xy"���&̠y�2�?2ᒠ��c.�b��  �rb$i��L$�� 7�4.OA5O@-O�~O#qO+no-{O* @ $Y� I'�� o$ޔ�$�u�ng�nh�k'Řn�&o�zVnp�&z� z�'И� �p�&lB"zoz�?Ż ��&z /�Ũn�&o.zoz�6z_"zpb{H.
�zzt�z'zzGzpb�lbA�&z/��t�z0����� p ���� � 6�� @o!ii�%i�=��(/`���iE ��bH
�!q����4"j�b��&�l6��"kjb�okm6�m���� �mD.E4nmb:5��c�o&o?"�nb�o ��p�l� � ���y����"� x��?� p%� � s�� @o�k �퀳� �i�l�&���j�魯����� ����O�e��U�lUI1w    �Ӹ U�T�@�	H��2ă���>��� @��@   x�/�w�!�⠵��!�T�/���a+�<��l��惠�x�lT�bw�c�Ʀ�l4�&�V΍�'�����/�$��Z$�$�wY ��h��<*$��R$�t��'����$�TRH
�*$� �RA&��+��l$$�wY  �H+)$��w��i+9,P���h,_���f��?�ˤĄB��̤���̄oC�����Vnw&��!��hw&��?���������$͕�+),�xl�D�2�� �  Sz ` �C\���� �(?���O�&,�-^���b(��(M�(�+����J,�������      ��&�
U�� y�r�b�g��w��~��~��~��~�Hr��b��l��fxf&2�&r�$&���Ѐ���$�s!i���!.q�/�D�4�&#�z-i�z��+� s�vOI `Lzd���#��%��z'�-�K()�E H
�*z�+���'�p�&#�Yl"z,i� ��� �$ݔ�� � ���ِ�r��"�/    �� `��d� ����D�فh�ٲ��K ��F���h�Ⲕ�K �����XH--sv /���^�(��a�/,-�W�/-(9��4(��@��-�?�$���6$�;��亀�-U2@��>H/�ê = L()� ���b
�ԉ��ً ��
.

�ٔ��-�� ��J�(�� ��I()��J� ��K�(K�(�� ��4�l.�?� �!�à����&,��!�㨊��4£�l�è���/�� �yd f �����C

�
��ɺ8ɱJ F (��Z(/�:�HG�K()�,�� � ���݁ls�Jts&3u&uuCH���u�u_��a�"��j J�����b=��D.��&�
.
:��3"ʁl�`0�����'��'��'��'�7�����r��{ ��3&�'�'� ��q�>��&��'��'��,�|�q⨙�貚�&����3&�&�ǎ�G��傾�� 	�&�H�	'��	'	>"	�dÁ�� ��������������������������<��D��IW�&�yOw��ˋ'��P\G>�U> �l�<�<� > ���r��s���$������q�!B�����|&�q�!>����|Xn||&�����'�����r��r�{����r��r��r��r��r��r��r��r��r��r��r��r��r��r��rրt�K�(՗����� ���<��3���ZY3�X�[Zf�Y�-�e,�k+�li�Eh�Ig�E��U�ᕒ<� �@@&Y�������'��'��'��'��'��'��'�����r��r��r��r�~�qr^�/�=�qKb(�                                                                                                      +ч^�"]�#r Uq�Yp�\��U��[��\p`Eo�Kn�L$/��������~��w�����r��r��r��r��r��|��'��'��'��'��'��'��'��'�����w��{ 7?^                                                                                        �o��U��U�I3,96 D˓3T�>V�UY ���r��r��|��'���q�/�������$I��������'��'��'��'��'��'��';�'��0��ɹ�`��K�(���p\? ���/���VQUISU                                                      ���6�D5��9�7MW���ǔY� U��^VE�K�L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���,$� )>��0� o%$���*$� )0�;o� ������m&�j��nb��b��ɠi�
���a��i�������7�Қ����b�����(��t�������� ����d������j�&�
&���֪
�J��z��3!��� � � ��� Yl�+ �Љ��@���� �A?ݹ�D �  ��& o�
c�ט�9��b�ט�/�e����(���4"�Vnn/��s��y
�6
�<��n

&^&O��H ���������װ�o>"
jb��i= @�&(?����9�ܘ  ���J� ��
���� ��4��l��6��C��d������|܊���� 怼�� ��"��/�c���� �(�6�� ������V��o"��i0��'�zĄp��¨������h z�p��¨�u�����h z�p����il'l?"
jb

r:
&m
'm�+ (���pF��6$ ���K ��b+N�(-� s�� �۠�#Ӛ��jz6� ���6��)���   ��K 	��
�� ����\�� �����k�y�(ώ��4�&Vn���S�'��ő�� ���i��b��/��� ����/���YH/��������龽b��&��"��bF�����b����D� �       UpHb�p�ƀ���k ���(�y�� ���b

�
X������bF�	��&� ��Pnl�(Y�lc@��lD�
�遬������������"�������c��c�S�	�#S�� ��ϋ���8��4� @��'��'$Ϟ����q������'��'��0Q�'��'�$���阶���$��������'��7��'�$�����7��7��7����C �DLN!M`�8��CA�	�	��RC! �Q 0�̓A�3�;�4� �������̉�Y����$�����q������'��'��0Q�'��'��7�$����������s��s�$y��顫���'��'�$�����r��r��{ ���r��r�{ 	��ߢ	'�	"�{	�"�{�����&��ھ��,��|�� p  ��BD�ާ%��(���s� �� &CS���3r%�,������H��Y�$Ƒ$��$��$�����P� �� ��  ����lXA�c�����X(C� S�R��D`���AŠ��c  ��DO�#�8(�#S�`C��E`V��� �N$ �U`���� �� @�΃�CA��S�E.1  �B2���T� E�`P��;Ʉ�8L`!�� ��P� �?$ ���48N�PӄMDQ���(���(/���(����t�����c���������(����/����Ѩ��(��(�����(��(��̏���� ���&!��"���� ����� ���(��(�Ѹ��&�􁀲��{����䂀���{�EfJ�n      $ ����������}�                                                                                                                                                                                                