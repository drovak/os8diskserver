����  � ? %##   %## ? %## %# ?  %#  %# ? %#  %#  	  .  %#  	.%## ? %## 	  ?  %#      %#                                                                                                                                                                                                 
 @� M�� ���    � H   � �<!
 DVD\dD � Cg����5�����                X$K ��#J�A             � ��  (�� ����������ϯ� �����	��@ ��?��� �� i�u�!��y�!����ϖ�r�� ��������ji`���j�bh*&*�6���gO�M�=��� ����.&���,��f!-�/,.�����Ϩ�����..�����ȟ��� �.-6..B*.d.,&*.6� �����-��� ��*6��C*�t� ���/1b00d�/��߫ ��/��K ��/��K ��/��K� K�3 ��.��&�.�.��b���� �����✜b���朏+��/ ���k    ���&�.e���+ �f(�!���c*�b*�t� � �I(�!��k���@��� �   ��c!��ˠO�ˤ�ײ� � 	h yz��x�d�/����J��   �4�����~�� � ���6�{I�����       ���6��C��d��6��N��7��D��J� �    ���6Ζd�>�̃�̄� �f�Π/�͢(�����ΣK��b(����/�Ͳ� ���/�G�<����"���H�*��"Hc�b�*      ����K �� �� �� !��� �"�� �&�� ��� ��� �%����K�������� |	G�m��|�G��|�G���|G����|G��� ���㟙d| ����m��|�����|��ԯߙ|���ݻ|���ݸ�� m	�|�G�ͯ|���ݯ��|G����|G����|��˸߶ �|5����|�����|��˸�� �|;����|�����|��˸�� �|A����|������ � �� �$��f�H/ 	��/�<)��J� � �<�� 	�o/㠎>i��"�� d�/�>��@�?� ��:����o:�?n@!l�"�9�j�ʷ ���@.?,  ��|�A���� ���4<ț ����Ϋ ��I�(��!�~Ș��J� �   �>���� ��>��|�A���� �yz����r�� �� �	��<� ����#��   ���I(�!�B�h��6�L8 ����C�e�����c��C����/�:K��㨶��?�>�@.? + �B�&�B�1�&��J��J� �   a�&�&#�����J���� .�1&116�������R�� � �>�c��i� �������m�m@����"�_#C� � �>�i������������ ��4捔6��I �� �m`�_�&��n٦<9��D���    �Ĩd��6��B�B�ń� .Ĺ� ���b�����Ź{      �����k      �������/�!� ��eb����+ ���r��r��r��{ ��� ����0����� #�#��"��" 	2` � ��8�� 	2�� �����!Ͼ	���Ͼ���	߾���߾!���)߾1���9߾I���Q�ʾ����� �ɾ&�?�� ���� 9&��9�/�!��"�9�k ��;i  ��mi;�  ���6� �� �4�i�4��� 2{��{Ɯ2�J�����2���K�  �Ip�v����~v��� ��p�v��uv����2�J�pv����p�~�v������ ����p�uv�������Lpu� ��������p� ���L ��2�J�DY�\qp� �o�������� pY�q� ���!"  ���&#UTo�����q�p�o��2�K��\qp� Ύ��qp�o�����qp��ʞ��'qY�q�p� ����qp�o�����q�p������q�po����d�ut�~v��s�v���~�v��2�J��ut�~ؚ�p�sݚ�s�~����^"���]&s~�v����~v������U��T��~�2�K��sv��������s�v�����D��sI~v������~�v��~~�~2��������� �� �����D� �p���� ������p �B�
� �2�J������� ����p� �2�J � � !.�/�� o�g���k�  �i�ys�~z��2�����ys�~z����6�ys�~u�z��z��2�J��ys�z~�����z����V2��ys�~z��y�sz��Ҫvƚ2�J��sy�~z��Ъ�s�Ӛ��csiu�y� ������2�wsiu� ��v ��2����T .KG��s�u��o���z�������o���2�������ʛ���o�������vɣ�� �qs�u����̰����o�����i��s�y~�uz��2����s�ɚ�2� ���ߘ�� y2 ���e�� ���b���8� �
2�K �ut�yz�xv�������� ����3	2�����s�v���x�  �2�����s�v���x�
������\s)v���w�!\� ��z���2����\s)v��w���sv��w���HǞ� X� ���y ��2�����y՚e�y~�z�2�J����yy�~z��z��2�����z������?�. ����2y~�z��yz����2�J���yz�������uyy� ��������yz��� ���| ��2�J��y�y�~z��2�������y2 x�Ji3�x���!J����x�  ��3��2������J���x���x������1 . � ���r � ��~z���2�J��r��r�~z����k��;z����q� ���o����4��q� ����o�2�J�z���<��q� μ��q���Ȃ�q�oΚ���W��q� ����q���ު��q�o��	���q��� ��~z����� ������o��2������ �����~z�����q��o���
���2 ���xJ�e�wz���D~izÚJ/��JJbe!D�/�2����w~��������˞� �5�2 y6�7ږz֚w8� �
2�J������ 	5�20y6�7��~�z�w8� �
2�J������ o�5�y6���37	�~iz��w8� �
3�J2�J��������"	��� =	m`��/{ל[<)�D�DOD�Ebb<E��G�<<�Z<)��U��Y/X�&mʚW/V�&{ߜ�D�{s�D�J{ ���{��m�UT"D{i�D��m�SR"D�bEEbFGb<<�b<)F�JZ<)DO�E�*� �!���� .!R
�4�{��m`��D&[<)H<)DOn����{���G���J���M���P���S	���V
���Y���\���_���b���e���h���k���n���q���t���w���z���}����������������� ��?�'�i������x ��
��
��
��
�� 
��!
��"'
m�|�����|�����4�i#�,����$:
{
�l���2��2���%F
k���2��2���&�m���2��2���'�
m�{��Q�)��&�2&��i 2���Jk�{����){��Q�&� � �<�/����r�k]"Ok$6�#   ��6�}I���(��!��b<)��Z`<)<<�Z<)��J�(��m�{��T�2{i|2ԡ��2�h���<�����<2���   ��6��B<�������)A y��D�b2�i�D�D2D�z�̀�>�i����������������Ϛ� {��۞���sGN"L   ���" �2Ί"��#� >��t��rq� y�{#�z��z��2�J��z���� y�{,�z��ws�v��d /���y{�Q{�2z٧w�J�iJa{_�Jd"�����A�j���B��� FG�JJ�NM�RP�VS�ZV�^Y�b\�f_�	jb�
ne�rh�vk�zn��q� �#�t��w��z��}������������������������5��6iy��P� 4�7��nz��w�CCb8 �����J���c���C/���������/� ��{�f��{ir���x�x�xd�/�4����������� �z�w��<����67�<����= "]O"�62 O*b
�ND�M�*b�ND��� *(��EEcLDE*t�С�������" 0��z�!v�!��"LDQSD � �� �� ߧ ۿ ÿ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ڰ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  � c?� c	�C��$�S%�?� c	�B�S�%�X?    �  ����  � /�?  I@��m�mm�@�/ ?p c	à��Tc���c��G�(R��5�cI���cӘ�@S�%�X?  c̘��cI���cØ�$�RS�cY���cט��4S�`RQ�5�cI���c˘B a�Tc?� c	SA�`@�e&���cC�(S cȐRC �T�E& �8`.A c	��@TX��4�TENn!c���c��ԀLUVBLN U�?@ c	   c�?  c�N%�XAR�ťD���c�	H�1:X?  `?P                                                                                                                                                                                                   