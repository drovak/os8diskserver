��� M �B ��                                       e7 ?< ?0?8=- =f P +���������                                                                                                                                                                                                                                                                                                          ���������������n��y��Ǡ������s(�����K��0�������?�������9����&��'��&��'�>����?����s��� �����'����Ι����ǚ��V���������� ���C(��c� �f2�U�����-�V��d�Hǥw���� B�N��K��\�FطHt��   ��c�(�������N�����"��������9��ǉ����0���������
>
����i��'��'�>�����Ǡ������{��<��|���� � ��c����l�H.�������|� � ��؃�惼� �    ����ǎ�����̦gWO`H�P ��\��t0���? ��������7��7��7��'��� ���������'��� ����@>�/��(�����!>�|����9� �
�����H��C �	�T� E��L S�ϟTI_� 0�ƟT���� 0����ƟL`!� 5�N �灼� �/1gK w�O��l߀���}���X��Yڮ	�֏  ���b��c��c���������2������I �
��"��c��'��"�����- P�!>��b(��J
�
�▧k ����ɐ�TX��C �	���N�`�a�4��&�����c�����"(���F.������� ��ş�R1��� 0��n&�����������0��o p�J� �/�0 ���?��������)�����b��c���[��0��������?�����������r��s��   ����r��c(���&�(?�˦�볻���?��������z    �������̟�O�#� 5�8�5 `   큞�� Wx�V����5�NT��V�h�`�N�������u��� �(����c���n����J
�
���c�����2P��������� ���"��c��'� � �	�����9��ǉ�Ɂ��!��������~�|��'�>����|����|��რ����<�|���ᴚ��4 ���C�VY�@���NdH��݀H�\��]��Wh�=E2AT_������ ����׀�

�
�耎8��J � (���� ��&���,�(/��������(��(�݄��(�׸��c�����t�����<���Ƞ/�����<�������n��r����+���� � �ݠ/�޲&!�Ӏ�� ���(��(� � ��T� ER���L���� � �=����	F�\N π��}��? �ҟC� ��h�8G   �n�b����0��/�����J����+   c�(/������������� ���bJ
�
��׿(� ���(����/�����GL*���OD�2���� � ������ ���� �����@� �t�@� ������?����0 @�/� �   ��c��(����/��D� �����ӓ���P�� ���?������������5TXL@!�ßN� R�3R�A� m�5C��1 ���i
@ `�Ƣ��{�ԟX��4� 5XS �Y���N$ �Q 0 ���� ���             �Ā��@�o�O 8pH���� ���������'��7��'��7��'��7��� ���������'��7��'��r��w��� �����r�r�r�r�|� ���l��'��'��'��'��'���                                    b�!P'   [���E��Z��c�F�˳�w�(�\_�\b�5��G�䬰����� ��  ��c��c��&��C��d�!>��l�������L� �  ��c��c��L�(/���(���(/���(����/����"��"��l�������*E MP TY                                                                         �����_E�\                                                                                                                                                                                                 ����ƀ�6��B��r(����o��'�F.����&�(?�����0��'��J    �	��)�����/�� � ����b����'�7��0 ������&�7�'D�'�7�7�'�'�'� ���
��޵�:�� ���K
 ��� 	 �Z����߫��
�[��@�� ���c�(/��D��&��)���ؠn��r���ـ������(����/�������Â���Ė*      ���ī+ ���� ���� �	������/�Ĳ� �   ���c���Ť��Ũ/퀸���� ���'������C� I�Z
��dTB�^��XNX9�� �\ �U���
�(���� ��� ���0��&�>��怀C�d��)���b��n��h����� � ���'��&� .��&��&�F.������/�<����Ð ������O������@��� ���������������/֝��������:��� ���O���8@��9����̚      �ê�H����������߀��\�� �   ����������� �������t� ������� �����(�
��7������ ������t�����/���� �� ������y D����
��K ���s� � Ί��'�!>��{����9���<�F.���� ���-��묀
  �      ��U?�܀�� ]�^��� p���E߼9 � ���Á�������)�
��'��z�8����� ������&��?�����b��c!���������D�����N��7�������̠      �����@���‐j  �������)���퐠���� ��޴�鳠��� �� �             ��U���ت�߫�B�����������E �� ���l�(?���J
���H!�扨ê����0�d��8����J
�

���J���    � ����/����>��ϻ�˨/������b�k Hˁ���t��K̀�� ���"�����'��9  ��ע��b!��� �  n��������� ����  �5��_W= P\E� ����� ����Y��)�����������9���� ���&��&��ǁ�����,��d��J��&��&�����y�i�l.�࿿7�B

����'��D�����'� � � ��� ����������6����)����9������8�����������G� ΋]��}��P  ��У �����\������� � ���/�������O��������4� ��������2(���(/��$�����+ ��� ���&� �  � �   � � ���Áΐ����2�����b��b

�
�ಮb���H?���� ���'ܨ?��� � �܁&��?��"��i��?��8�� ��2�����]�E ��?���ߣ�� ��� ���6��B��bl��C�
�

�����L��<�����D�����|��<���>��だπ�����&��'��B��t��'� �� �� ��+    ����������J
�����b(��@������ˋ�ˋ��   ��� �틜�� ��
.
B�,x�VUG�M���� �?� �� � ����                                                                                                 ���/��������y����F>�����0�|�<��w�|�<��s�ꛋ������ FHGZ��\��M�^���׋N��� �� ���̀����9�
��Á�ϝ���������8������y �����۩ D���� ���<(����b��b
����.����� ��(����b��b��t»J� �      ��b��b�H/�Ĥ����b��t��'��K��ˀ � �� ����}�� ]5���_�:�0�F  �K�	��E �X��  ΁\�                                                                                                                                                                                                