����  �. #30:   ,    /	.                                                                                           
: *  
 *  	/>/=                                                                                                                                                                                                 
 alwo y                ? @� �   (���������}n�PH�������������߀YEZ�yw\�k�`����"�&*�.2�6:�?D�IN�RV�Zڈ��ag"ms"y;!�⣀�̎��ـȆ���������                                       P� ��f��H��U�3���f��A�U	5����f�iA�U7����Q��f�i%�� `�U�9����fMiAU�;��q�/f&MB�<�C�U=����f�i'�� `�U�?���f�M��;I�@U�A��R��Z �   @a�^�rU)C���/����Z �    ]	a�^r�UE����SԚ� � ,
 s��i��k&i"iMii<)� �k�J� ��i6��Cj�div6Mv�� �ijD��� H	FE�GL�KI�<=�> �  $  h  �  F���  gfb!g����V'�z���������V'��7�6'��)�PI��M�����窤Ԭ�� �AP�CrR�	1G                              X	x�� � @]_�`c��e� a	 e)^	 _�d�` �c �]r�UG���UI���@UiK���U�M��Q���@�UO���UQ��R���US���UU��S���UW��Z�T� @]a� ^I_I�`e�a	 e) a	 dI`	 ^�a �]r�UY��T��W�� �&B"� �P? ?`��؇��� � ���dX|����   ]	_`�c��e �a �e�c �e�^ �_d�`	 c� ]	r�+ Z	�� @]_�`e�c	�e�a	 ])^_�d�` �c��r�+ Z	�� @]_�`e� a	 e)c	 d	^	 _�d�` �c �]r�� ������ ������ ������� ������ ������� W	�i&��X ����   @e�_	 a�]	�h&rU)[����Z �� �@X� ��� � @e�_ �b�a��rU)]����iO����Q��W��i&�Xi ��� � @e�_ �a��]ŒhrbU_����Z� � @X ����   @eI_	 b�a	�� 3���o �4i)3�&���2�r�� 71�rU)a����iO����R��W���6� ���"��"�  WZ��� @y]i_`�e�` �c��]a�@r�Uc��W�Z �� �@y�WZ� �� @yei^	 a�@]�c��rU)e��WZ� � @yXi �� � @Z �� �@y�e�^ �a@�]c��r�Ug��W�Q����� �
��)��&�@���E��� 0�H> W	X ����� �@]�e�c �d�_ �d�` �]r�Ui��W�X ����� �@Z�  � @e�` �a �]c�rUk��Q��W�i&X ����� �@i��Z�    @yZi��� @yei`	 ^�c��a �a@�rU)m��R��W�� Z	    @�u�H��M����� �v �J
�
��(��H��� W	q�/�[� �� @a�]r�Uo��W��,����Z �� �@]� a	rUq��޹WZ� � @;]�a�rU)s��Q���@�Uu��٨�@�Uw��٨� ���6��Iy�O�Xi �����  y\i d	a	r�� ��ٛW+,wX ����� �@e�`	 b�a	 r�Uy��R�����@L@@F����2W��+Xy ���� @WX� ����� @e�` �c �a �rU){��WX� ����� @e�` �c��a �rU)}��WX�  ���� @:*��+��K�e�` �a�rU)��S��� �U���ݨ�U����TʚW���k   ��6� .�WiY ���� @W�Y ���� @ei`	 a�r���KuET �@@�U���Ȩ@@�U�����@@�U���Q��Ȩ@@DU���Ȩ@@HU���R����@@JU���S��W�� ���6��C��dWX� �����  y\i e	`	 ]�a@�r�+ ���d��6�WIX ����� �  \ �c��e�c �d�^ �d�` �]r�� ��!l��{�/�{��&,���   ���7���� �WX� ����� @ \�@e�_	 a� d)`	 ]�rU)���Q���X� ����� @ \�@e�^	 ]�a@�rU)���R���X� ����� @ \�@dI_	 c� ]	rU)���S��W�� W	���X ����� �@ބ�Ы   �����d�9������� �(����#"���5��""���"7�    �� �Q��� � R	���� �S����� T��W�� ����h�c��d�D>�/ k��Bi�bjjd�j'jkBjiti�JWY� ֏� �@e�^ �]r�U������i&�j&j�B j�jkB j�iiD�W�Y ����UQ@eI^	 ]�rU)��ڀ��i�bxxd�f&x�8xkBfxc�i�i�J� �U�� �� ���� q���W�i�f�h&��bH� O������"��b��h�k&� ��k��Ԩ׫�r�Yy �� �@[ ���@Y� �� ��G���U9����W�����i$��� �H�����h<��k ��D!��Դ6��K��������������� �� �ut�yz�xv�������� ����3 q�����U������U��ڻ���U���Q��W��-砟�Y������@W�Y � � @eI`	 c�rU���R��W�� ���6W[�  � @
yei`	 ]�a@�r�$� �����[i  � @e�` �a �r�$� �F������� � �� ���b ����+ �
��?�. �� 0	_��#W�X ����� �@Z��   @]a� aI ]^e� a	 rU�� ��cP��vf�H�� U驨�Z �   a�r�U���Z�  �  a�rU)���Z �� � air�U���W��#�X � �� �@:�AH��*��+��נU���� �#W� ������d0 ��� �k�M����   0Þ�:�fo�{�?U���ڍ� ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ��޸ ����� �ҿۿ�K ��Ĵ� ������K ��޸ ��޸ ��޸ ��޸ x�"�n�g&gg6��6g�&V+��P��x��x� �
� �             E	������ G	������ F	������ H	������ A	�!��4���� �C��!�㣠O���� ?	!����议K ���(�n ��r�rtbo�/�M�pt� �� �t�&��$��D��       �{�/�!���{lJ>����ul� ��u�� ��I����u�k s<r�!t&� � ��n�n("�|��'��'��'/o�|�n{o�0�����j~|f�}��!b��b��b�b~b��b����DOƄ����2�0.���6��6넟��������J�J�o��ߤ�2)�3s�0y>4�0�3��{}f1�� ����       1   BA�� � O�E�*� �!���� .!��zof0N���i=��,��;��< �7��-9� �}�/���s�� 5	���|�k�.��?���� ��!�!��P���J��b�D!����&�s��,�� ��z��=��,��;�� �s<)A����0X��M�5�������i,��s��(�� ��j�(�� ���� D����� ���+ 	 ��F�J���s� ��&�� �D��hF� �(�&��h
 ��O�D��摷����/2��3s�0yP��s5�v-� 7������&�5�� � �=
 �	!�o�k��QR�0D�Ƀ� ����b$�/8��%"��9��7����/�ʣ(��@����/����ʤ��J���&�/���'�/�ʤ��6� � �`k�6�# ��6'��6��?���M���PI�|�����>����|F��K0F�4���}�1 ������(����k ��92��9��r2�3�7� B�!b��b��b�Xn�o�Ϡ�����b������6�����X���d��J��'0��� ���ݸ л��   � �    � ����R����q?� ����� &1���	� f��� �g�(� h��� �?֘כ @	�C�� �B֘C�; C	�Ƅ� �A֘ͯK D	ք�� �x�(�� v�I�� �w�(��� � �& ��c��c� ���K ���6��0��7��C����t�2)�3c��t��'��B��t��   :� zn�����?�lnm�l� 6/!��"��{����$(/8��(9��(/���(����/�u����1����� �gVi)��m.l,  � ���&��&��&��D��6��7պJ� ������b��b��d��C��c��t�ë� �    �                        �w�kxU��U��UEZ�[\�]*�akw�]O"�62 0	��Ħ0�������q�ji�"��� q��"J
�ns&�2)ü'q�/�"�0y#�� ��iib7i�� ��&�ȯ�i'"���i ��K(*��I�G2�' �   ��bΘ��b�ŋ �� ��b�����+      0���}� f&pg&��'�U'�/� ���My0��1T��k�L ��7��77���� ���(���� ���⚬�ÿ� ���(��� ���(ÿ� pp&�6�F��s�<˘H��M�:�� ;@����7��4��{ s�<�� �=9 �9s <�� ��f�A�(��U-� ��f�k   ��"�hFޚI�:����D��� E	��F�y.�y�Eꛐ��pg&V1� M��0�V}�MW�1>�C�� �%*�/4�9�����3  E� V� g� p����������������A��B�C��D�~E3�A�B C0D0E�F0G0H�<I J0�0~�0~�0~�0~�0~�0~�0~�0~�0~�0~�4��4��4��4�1~1~1~A1~B1~C1~�1�1���1�1�1�1\�1\�1�1�1�1�1�1�1\�1\�1222A2�B2�C6��6��2~�2~�2~�2~3~3~3~3~3~3~3~ 0    �                                                                                                     �x�`���4 5�HR ���I�Cp-��Pc  ĉ���_ ���`�C� ӈTP��(��5��(�S�  P�ӈLC Q�T�A��8�S�� @   � �ぁ SR�� @� �  �   � p� p�ԃ ��!�Ԉ�z� ��L@8� ���X�N`!TԀ;����TX�	3� ;�8CUn 0����zM��`1�TR`�SB�HTX�	3�8T "��PM�[������D�8�AV`!�R@X�O3� [A�3LT�	 �Ơ1	�3�Ը�����4 B�4P���D��H��@A�ϔNE%� �                                                                  ��&��� ���b� ���fo�&o�c��d��6��C��d   �t�t�c!�⨲���J��J�o&ot"���Mp�t N� � ��;�=?�@<�>C�DF�GH�EB�IM�LK�PN�J���������ę�ʙ����H�49 ;B DF ါ         ((�  pp�pp�pp�p(�$  >                                                                                                                                                                                                