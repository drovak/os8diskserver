��� L @A >/859
8
8
9	4	3/W3> 2  0?8 **?  :2X   : 2?2>"""=> *	!!#<8!#;2
':   /9  .   82? 28*+/9++887			8
8
87
		6)                                                                                                                                                                                                �֔ D�h�P.������cf�s��s�������!���0��'��P��Á@λ��J�Z��'��'����@������ �b

�
��b����	� "�k ��b���Ϋ�J��&=Oy��@r)������j0"03d�Ҫ���� �?  �e��ǀ��`8�у\��E�  ���&��6��0�����D��J��˶ .D���n��&�T.��j��7��ⷠn��&��J��2��s��'����b��~��7� �    ������bŉlV�<�*��~��V�<�U�   �
��r�h���V�0���VT0V�z��F�����sP����ŀ��`�~����&��\�~� �_�W  c �W��� ���6��C��d��6��L��&�� �����   ��l�
�    ���&�����c��c��c��c�(��&��0��'��<���  ���Él��<���   �
��'��'��'��'��'��'� � �         ��D����� �(/���X�&��U�I��Lf a� c�mXe�������������� ����l��&��<(������ ���L��<ҡd��N��b�� `� � ����ǁl��������&�F>�����J��C��
��D�����J
�����4�  � �    ���ɀ� ������ J
�
I���&��&��&�ٲV ��b��b��k��O���~ �&�π���� ] ^�^������ ����l��(����� �����"��h�!>�&��<��X P� �� ��������l��˫*�ƺ������7��B

�����'��B��d�� �D���oɩt� �       ��� (��J
�
I��@n��#����� �� `�̲��&��&��&� �l�� ��D�W� ��\�W�C?P��                                                                                                                                                                                                