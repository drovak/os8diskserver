��� �D C �@                                                                                                                                      
                                                                                                                                                                                                                               ������G����&��0�������?嘊ߨ?�����0�d��0��d��6�B���������/���䖔�DV�	��� 5��CU� A����?���� �����c��b� �f������K��0���D� �         �N��{������ �T�G� ���V��`�d�����@ ���d��(�����(���   

�
�� � (���� ��)��K ���6��B�����(� ��(��������霋 ���/������(� �   &!����� ����(/�����������(��(��B���� ����σDA� �� ���)��)� ���(��(������ �   �� ޅ���?  ������i��J��9� � ������&��?����������9��c(��v�(?��'��9� ���'� /�&� ���&��&��@V�{&��'���T� ER���I� ��!.�6@.�/���"�k ���   ��0`B�D��F@�o��V�?��FGG��`�����P � ��˅�W��&��˶�r��j��bF�����rJ
��බ7��D��D��&��J�������ô�i� � ���T���         ��?�� �            �É�� ���9��C�̛   "@��� �                                ?�yc�FIU�V0�U ����P ��/����/��������c(���d�&b�&����J� � ���c(���d��4�ib!�����)������(���H����� ��f� �(���H/��@������"À���)� �T5Ӌ��D� P �	mm� �	��� ��㴀�H����? ��G�Su�@P�V���P�ϟTT Q��Q 0����T� E�S(A-�3 ��ԟX��4� 5XS �[ ���r��r��r��{ ���d��6��C��d���    �
���ɐ�TX��C � ��b��o� �                                                ���U�U� U��_B�D ����b��f�(?�@��/�����j���(/����؞��d���D�������       ��
.��б(� ������ ���)������   ��b���ɾ��ɘ� ��/��) � ���'��'��'��É�¨����+�N��8Se`1��P � .�H�-�) 6�����@�0� �����2(����&��6��)�� ���)��)���   ��&�� U@d�D �@��D�A��  �@ �S3 QP�4@S �D������A��B��C�ā�Ă�ă������Ø�p  �/�����������Nԓ�Se`2D  � �            .TF�Pb P�D��P�?y  �(����b��&��2����.��b��&��"��i�� ���/���H�6��/����� 0�������� ��&��i�i���?������)�9�/���/���虠���������9��DD�J䀛��J�Iƺ���Ř (g������y� ��
�� � s`0@Qct ����/�����M`Tă`���`��"�8��8ŀD���M�`HŀD��� ��&��?��"�c�&�&�&� � ���)��)��)� �
>�໻bF���i(O�����K����K�B�D�T2� 0� �    .(bu?�u ?@�6��P���� dD����DB������扬��6��C��b�D����b���� J
�����"��bJ����b�J!���b�?��!���.��b���.��b���Ͼ;�ѓ��&��6��0J��>�ςl��y  ����� c ���B��w�H.�   ���b��l�(?����2������ � �ڇ�xf	����Hb��Z�?�s �    
                               ��I��
��I�/��I� 
��I��
��I���I�/
��I�'
��I� 
��I�&                    	                                                      @V 	
�D 9
 D 9
� @
5 I
� NP:�8Lˆ8L��8LK�8L����������8\�	�3�^   ^�ځ    �NP:�3   �N ��1L�
^ �
�r\   �1L���2L$ ��pP��            P                                                                                                                                                                                                          �	�/�����hA�☙�� ���"��� ���<�����*�0��&�@>��/��:   �!�@����� �����c��Ҁ>�׀>����	��J� ������t����C�ś                                                         ��� �u �� �b ���(����n�J.
��&��"�������)��"��e�����D�k �	�/����b

�
�� ����)��)��� �                                                                                           b�T��U�u(p �                                                                                                                                                                                                                                                                                                                                                                                                 ���b�
�����������H�k �������� �&�É�� ���	�b��l	�<b۸�����J��� � ���b�������(�(/�������������(�������(/�鲨��� �                  ����V� ��k}D���h?��	�<�/�!��&��0�'
>��.�k���c���~�0����nD.&���
.��� �                                                                                                               ��
��� 
���������D���)ˢ� �	�/���(��k� � ����2�@2����6C5� � S���1��5���=H@=Ȁ=��=� �  @�����H/��"�˛�2���� �                                          y�0��bU�#[                                                                                                                                                                                                 �	  8�	�/�����f��f��n��d�̆�͆�ΆЀ��φ��&Ш��Ϣ!����&�(��!���&ɳJ�!���&��D�΢���� .Π/����� ��*������                �։<��K                                                   � � �� �� ����(?�P����L�S	� 0�P>��������㨪���ɇC ��P����GE��4���P�����`A���  �/���H�����( ��P>���P�	SQ@����?΀� �	�!>P�����d	����5��K                                     O
JH��KJG�� Iz ���y@�␛��(�����������(����@�☛��蟀���D�R�C� @� � ���bg��J� ���&��bc�����J���EVC`���4 ����� ��`A����$��4 ���� �(���כ���� 0� �                         (�H��_C��  � ��PV�                                                                                                                                                                                                