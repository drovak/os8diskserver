���  � �"=&=*=.  {/< "" 8 +?+8+*% 8??| < ??   <??   <??0   <??   <??   <.??   </??   >??   <>?>     <???0   =??   =?=   0   =??   =?=   0   =.??   =/??                                                                                                                                                                                                 �+&@ �� �����[O.y P �                   ������                           O � �8ƻe�b��&���� �p�O�m��B� �TO2�*;�� � -���w� a            � �����s�
��� �v���? ���?���R��` |B)�;�2f&&�&6&�&�&���t���;������� .�&�&%/�?�2�>Z�\+&],&8�$'%B�|�/����&A�@��Bi�����D���� ?�Ҫk<X�E��Kß�E����&�?d��F��;����@�����  ;���{0 c�s�9�!6���Ā���[�<��XE�HI�.�/�>�Z.����@)�/"@K��G��X�>Z�.��J���"�<��E�2Bi���(����/���@E����E�?GU�A=�Z�j��&EH�P.����;��HK������*D=�qк��*DE�HP�X.�F��@��2�/G�@G�<����� �2�/�\��@)]@)� �   �
P�@�� @+ 	_�IdL��.������&M������X�Ni����K��������&N���0(��@���Xn!.7�Bt'�K��G�� ��/���@.��/�;�	HL�N����>���/�R�Ri�Ri�@)�7�@��F�@)d�@�X$�t%'��6Zi!.7�/G;��H;  \ t��8���  ��XI�F��\Xi�\�!���XI�!���t�&f�Kܟ�X�.Kiة�L��D.�����$�;�DH[$�����"H��Q)M�����"!2���4\�ipO�x�_28(�|R8�2t�.��|KԟG���rL���v'�+� D. b ��l�Ub!�l!t=��!�z�<"�i;)�f��H/ZL���1f.���>��&L��hࠫ�N�Q�Q�Q1�M�����\1b!���i O	x�_�;�H
&1"�&8X�r2d�9��9b�9r�F�@)2@)0&1 .1b!1�1�*�R�b�R��R��l'"
��JX�
X~$
'%
'��0bKië�EH�P��k �88�0�uO6�<�|1D���@�X$�22t%2'��bZiGV�����K��G��W�G\�x�\b!\� �� ��6�B))&�"��i �9�l.��t9�'8��r�l88t���&9�&�|�v�<X�EH�I.�>.�����@)Z.���J���/"@K��G�� �F u�u 0  ��Q��[��Dx�<L������N�7Ki����&�&D�B���A�=������=i��J�ܖ�@)�2&B��ݲ�b�i�x���6X�$'%'X����@)�� F2�@�@ے@7��@)7Q)�Q)�Q)Q)BZi6&H����b� �    ����� �@��@L������;U�Z�N�@H�`� 8���F���f<E�HB��F��Bi���bc(���c�/�E�H��&�?���FA�=ߓ�?����@)@)GD�=����;F�H��F>��U�(?�ɦ2����<������&� �2Ki���EH�2�/�K����P.��;���3�b@ɛ3�/���@3��?��>����<?��>��"@�@G�;��H �A� v��`X ��d��4��b98h��6��C��b(����	&��&�	�a���?�䤘��ƛ9&��K����&�9&�d���"��h ��Ǜ'8���~��&���r9�b	�l	�<�tǁ�� �a.���ϘO϶���&��&�d�;��K       ����(���/���歿���� �����x[� \F\�D\�]\&F.�� `��)3U).U)NU)�R��b\&��@����,��<b�|��[�������&�\"�����b�l(?�!�\$���D�J�!�l�\�t��*��&��*<���Ki���KI�����D�E�HP�.�/�;���@G�,<�L\�    ttIdj�T# Z"@! �I�   Q)&�Q)Q�Ȥ�B��(/��� ���Q)������E��Kן��;P��U�L��N�Ti��� ��S�S��B���� ��B����/�(/U���bc(��c�/�R�(��c!����Q)Q)��F͚U�FR� ��R�Rik;O�� � ��(0 o�'�*4 � �^Rf�������T���Q�Q�Q�R�QE��I�Z.ਢ�JT��.�>��/@)[-"DM͚�R�RiRiRib����J
��l�0 ��#�z!�����S)S)T�����&;ӔR���R�Rik�������/�V��O�r�_�ǚW��\.x��Ot� �	X��  ��x����� �f� ��/���;��� �Ti���\Oix�_���/�P�8���X.��/�Z���.�>h��@��8�.6��.�/�>�\@/È�@[�.'X~.-�Z�9� F��@��� E	�P�.�/�;��H ����@)�+ �3�k<�����@G� �@R�7�kJ��@�����	�I� �8 R�e `?����&�6�6>)d�bc�c��b��[ ���Z�ਥ�J���H.[ �����2@��Z�.��J���C/@)X.���/��.�/�[�'�{��2�;�T�;6 �d�b		c.	c/.b��T��P��f��*Vn�b�iɀ�       <	>����"@G�!����>�� B	���@���H/�����KU�� B	���@������KU�� Y��]]bD�⺚d�&\Yi�^��_&]D.]\b\�_�J]^"]d�O� ��X� ���&8�'�9��F�k8�rg�;�D�; � �H/��"�؋ �!��&����<E�HP�.�/;���@)G � ߠ�8�Z
P�?�� �&���k ����k�C� ��&�&� ��&�&� ��J����(/�����K ��n&��; �"Ȳ�;� ��r�/��� B	���(�� ��(���U�� �I.�>.�[��Z�.��J���"/@)���
D
�
C
�
�  ���� �       �I������ � ���\FOn������\FOp����� � �"b8�� ē�� !�&8(�|!�K� ��2��F�[0���X����s���>��@)�$��{  � �d������Ë����Ë;Ӕ� �dn&	&	H?�[�����/��"	@9���@)� �  Ӏ �e�K e��(� �� ��  ��A \]f^_f�dbeBi��� Y����i]Ba^bb_bc�i����a�b�bc�i�����B����/���U��/�B��������Bi��� �	��/��!�U��\&����!�@��!���*�b��b	b(��H���	`6	a6	b6	c6�ך	�"֌������K ������Ȟ�# ��O���$� ������������0��&��<����t��D�����c��ǉ�Á�ǉ�ĸ�D��J��,��r��|��ɻ�"�����'��'���8��: ���� ���ɮ풌�Ɓ���(�J�����F���� `� >��b�8p� ?��"�����'��J������ ��.��qߧ�W> nb����8� D���� ��Á������&��Á�π��D������c����lЉ<�t���	�(����n���   ��.�ǁ�ʁ����r 𿺢���|�����v ��Ʋ��r&�b��{� ��&�&&�J
�
���9D�����!��ѫ�� �E`  �����h�F�=V�8������ \``&]�&^�&��&]^f_�i�H.��b������J`\&���    ](^�(_���]� ��^(/_�/Ȟ����\\&�\�� ���&f��@��q>ǰ~��&��J� � �	`!.\`&��&].�a������(띂��.��i��J`\&�]&�^&_�h� �@c�__&b�^^&a�]]&� ��@_� Y��cbDD�D.c�* ]H]�^.^_b_�\�K� �_D._^b^�].]�k �(�� ��U�� �Kޟ���\�b�b�h�F���x��t�JBɚ��/�;�S�K�2�{ C	ɯ� ��CЛ��/�U�����\��K -���-�/��"@X�--&� ��߲��� � q��?�"  �]�� X��\Yi��]Bi��� ��X�Bi�����/Z(�U��d�A�\F.�]Xi�]�]Xi�^�]�"����&(?�]����^2���6�&���JD��^�* ����J
�
����9��B���+�(,�(��)��)� �]fn]bF�]]b�� ����?������ݫ `-�0�� ��p� r8r����    @   �   � �6p���k��A-�Pʪ�#L�SS5u���g�u�o�_��_�֏��_�o�?  � ����� ��������8��1������/���.����N���?����^���O�r���;��_�9�n7��~�/,��o��������    �    - � =   M � ]   m � }   � � �   � � �   � � �   � � � ����ҷ������C�O� �����������Ĺ����g��������l�������� ������!����������?�����/����R�������V�?��������������`��������q�������u�������������t��������o����������� ���������    � �%O$ N��J�����b��b��ǁ�Ħ ����   ½�ƹK;Ɠ � �q�8x �T����Zn����D!���b�&
&PX�.[w
7��J��;   B���(?�OU���F ����� � �ۮJڠ/�ݢA��o��I�� �
��Bۃb��bށj���;E���'��'��Á(�����@�   ���������c�J
��

���J��0��d��0(���(/���(���(/��(���(/��(����$� � �      ��4��c@���B����O�߫ �� B� ��o�����χ������<�����������l(?�&��<�&r��|�<��z��Á�����֚��'������<��Z
��|�<��|�(6�*6�<�&|ܾJ��J�
&�	&�X�
	t��	
g	�J�����r��{&;��!L�� � � �$� 3X���������������������=�FڋA��@ � ���0(��H
��桁��.�ࡐ&��� ���'8� ��ݠ/�����t������''b!�� '⠶���'��'��'��'��'����\Zn]Oir�_����b
�c�(OH
�f����b���4
t�O�x P� �� �Z^b�fj�n �    O ��D���[ ����� P��?�ø������8� ��  @��  @��  ���  @��  H.��  @/��  H���  @>��   ?� � N� � O� �  � ^� � _� �  L n�� � o� � ~�� � � � �� � �� �   ������ �D�� �� ����F �����������F���O�� ��=�                                                                                                                                                                                                