��� L �@ ��/  m2> . ) *+< ?)? )) ?2n 7���������                                                                                                                                                                                                                                                                                                                                   ����C �\��0�L�����&G6��cHc@@b
���J@b����w�����r�@rJ
���!E�K�k ���&��6��0�����D�J���� .D����n��&�T.��j��7����n��&��J��2��s��'�����b�~��7� �    ��    5���>���
����p� �� �L�/��"F�b������BKbHI&J�)���C�b������K�<I�b����ĘK NC�JL�/�B���BO�������B��E���F�J��)����G��������� �@IbD�I�I� ��)I@$ɀ��Ѹ	
&
�"-b��

r!	⠛���ʏ&)O&)������I��L���� �
�J�@����� ���6��C��d��6��L��&�� �����   ��l�
�    ���&�����c��c��c��c�(��&��0��'��<���  ���Él��<���   �
��'��'��'��'��'��'� � �         ��D����� ���D	�c�怺���I��La��c�mX��������������� ����l��&��<(������ ���L��<ҡd��N��b�� `� � ����ǁl��������&�F>�����J��C��
��D�����J
�����4�  � �    ���ɀ� ������ J
�
I���&��&��&�³��d��l� �    �~�(���������� ] ��^������ ����l��(����� �����"��h�!>�&��<��X �� �� ��������l��˫*�ƺ������7��B

�����'��B��d�� �D���oɩt� �       ��� (��J
�
I��@n��#����퀘� ��̲��&��&��&� ���K ����D��� ��\
�W�C?���                                                                                                                                                                                                