����  @ �� ��    	  	     	     /           	/      :     :     =      g;            n  u8                  A<?( 	���������                                                                                                                                                                                                         	� �@ٔ�MA    ! � ��       D�x2� �         �        �3   � �� �          �	  �  �7%} �               �6��4    ����dB� ��(�?��s�@: ��M��8m�e��a��$���g2�� ��`���f�M(� ����,+&&����/�*��)�!����:� &�����ÁJ���L���/�b/bGbH bHHt.E&�������c���F����F /�cF�c ��@6�D6�C6�F�����F&DT.F�@���F��i� � �v�� �� �� �� �A]  ��|��خ� ����������� E �� ����D�/�G�HED�������<GGsHGtHED��� �	
�&l&�+ 4��4,��� ��&&b� �4�h!4�&�ί ���6��B��  �
��� ��� �����)��)!��֫���s�5t�9�e�h2��c��z�!.�/�/�b����naih �   �/�}��*�/����r�;&�N6<���/bF.bEcFFtE�JC�8b����M)@�(/���鴢?f!.��iA>#�#i��� (?�D���M"�<����/�Ҩ�8��"�L��L����)<�ҭ� ��b�E&E�6L ���);��<�����J( � �K/�JL��N�K"��?����� @��A	="�/�?���N*b����O&��M8����@��/�L��"�E&EA"�EbHr!H�HHtH8r �*�/���),�!+⠶��Έ#��� �(���>��J�/�"�+�J�*��)�L���� �E:bO�E�Jά� �OΘ�Έ,+&؀���B(��X')��� X"'ӛ�t�O\�'e�'� Y��` 0/�A�� ;	(���(/�H�����&"����k�ꖦ��;�!⠐�;!��/��ȏ���J *��6.b��n�;i!!t&)�J�!�!�h�J;�&!.6�/ɠ���bȏ��&�77t� �!F>�!!CJ
����� >s���!!4s�!��K    � W	V��7 /W\�(7��� Q��� ����O���JO)O)� ��!&�7&&f�&� ����� 6.�&�8J>
���� ��b����bOВ��8�0J
��
.
O�4)�0O4��΢J6O)6)��      E�bFEb
H��F�J$��6.6�kL� �� �� �� Š  /��xR()\()0a./�/� ���� ��N �E�dE
>

�E�8�E�� ��(����H/��"��� �������LÙ" �GGbE�nFEc

�
��E����EFD�ŢGE&E�?�¢�E�

�
��E����)� �E�.F&E.E�G�E� ��)GH.F�J��)�۲   |r zw yz xw || ~| zt sy oy �� �� � �/�@ �?� 8���.E&*�/�/bFc!F㠨�FED�?�!>㨀�Lʙ?�)Lϙ>�9��)<����Lʙ/J)Lϙ.J�� E�F&E !D�E"JH��F�JH��Fb�F�.�F� F� !D�"FbJ
�bHH�FFb!D�F&���ց<$���;�/A��!@�������}R��_��0��� �c����E&C���E�J�-� ��/b�b�Nb���N9 : �   ���A�b�kL����)NK)/J)"�1/b0   ��%
��NB��A��CF�P��7��`����7Qx��7�[�ur��h��/�ⲲP��_"���e�*��~,�(/��lr����$t	c%� �)����ɥ��%�� 6�G� �@�����G���� E�	&�6��CF�d�H6��CG�l ?E�L	rH&G�JE�/�F�	�b�cEc		wE�J	�t� ��E6�@N�@ C�/�E�(��F�nFEtEE4(��GGcE!E�?F�z̥&@��tO��t���( L"�|���� ���g{�������j �)|������ ���_�ص�7� ���n� ��i��6��C����90F���"��d��6# �  @������LÙ��EEcK/����/J)��)��/������ � �/���?�J�''�'}������~ /�ӂ�*���
� �    <bR��b��&�M"F�I���&�P.��/�󩀀�ۈ/���H���!&�H+�E&y/�� 6 9 FFb�E&�EÁ Ϙ�F�/��"�Fb�:�  ���#�kL����)" �9�EEc�Li �tq�5d�b�o�bl!l ���s�b��bk�he�2b�� �"(����/�ؾ�|�2�J&c�bbb�j!.�/�b�d����w����w�p��fـfɔbFCq�T�ɓ��/=/��N6N�&�'&/�?���MA��'c�l��<�h" ����"����y��j�������&�	&��&��!	㠸��J����D��������K���K����/"粠����"��E�lE�<�	�E�lE�<�����ڮ�"{             �b�c�� �k�h�PH� � ����5 �U��HA��90N/c���N�"EEcAf���M;��6�!Nb1n2�i�������&C!�⠞��6���7�t��u��p<�t���A@�� p7 p��)�� ?�!������)$�/��������;��6����}����bz�.o ���m &#6#\� .W �b�i��k���Db�`�� �/1�'� x�p�A� �/��&d&�"����&B� �����F�E�h���EE&���������E�$� �G&����F�����E&E� ���G&�F�F�E�*�FB� ����k E@�E�/����E�??bA3&�1�($��k �?�(� �$�/���1(�!�?.�$�� �$�/"��1("���
�t�����7W�P�?T ,0�b~i}&&b�(/���(|��(/��� ����)��)����/�,�!0⨅��0�0�n&��)�&��&���/�&�t0�J�!>�bi� ��ƚ������.� ��� �����)����� ��#E�lE�<� �Eb�F6E�,F�|�$�㜵����p�`ܖ�/����v�� �	;���6b��f;6 !样��6��/��� ����&��/����/�����/�?������f�)���/������� �   �	&�F.����l� ��/�	�	c	c	c�l� �                                                   ~ �U; �7�QɃ��p[��PP3   ����    \	`d�hl�pt�x|����������������@ �  *@   8C    �@  �@                                                        ��D   �   zV   :5   p� �q� �r� �s� �t� �u� �v� �w� �:D   �D   ĺ   N �8P`   N��C h SσG�҃  ��DX��C  �/ 5R�� @ S� @ o�R1��D   �D1� � �N:Q  �� B�      ����#�##s�%&�%'�!.%�"�S���b��f��&C &~�*7�xqO�         ��tiq ���/���t��|+�!��+�+b���+�"��� �"(����/�� +�+ `|����"�tig�����e��/�b�p�� b	c ���|�� /��	r	r	r	�|�H�#�n&�"���#'���k�H+� b�@.��/��K�E	�g����� �"@������%
�F������	�D�                                                                                                                                                                                                tq�)(/��8�7b�^r(��v)}��#&#-"-#b'�}'	#�!.b@���#�J�#��縲q�&`{�/�����q�!�&���"5f�!�)�/� ���|ɚ���Y��Zb
�j��J���� �
�~|i �/�]�)��!�t �G�/� ����� ���K��� �   v*&��p��"          	  	     	     /           	/      :     :     =      g;            n  u8                  A<?( 	���������         ��Ž���������Խ�������ӽ���������ƽ���������ý���������½���������ƽ������������ӽ����������̽����������ؽ���������Ϲ�������������ω����ŉ���������ӽӰ��ĭӰ��Ǎ�������������������             �
����Ͻ������������̠������̍�����˽������������̠��̠��ҍ������˽��������̠��̠������ҍ������Ƚ���������н��������ҽ��������Ž���������Ž���������Ž��������ҽ��������ν����������Խ���������