����  8  0  (       � � �    @   ��&��� ������è�/���ҫ���h� ���������� 𗭢��h� �� � ��(�������J#���6��Cвd��6��Cϲd��6��LЉ<��t �� ��É����    ���bЁl��2@������0��'��J                                                                                                                                                                                                � ;�2��E�uUE5��E ]�* a!. �^Q'. ]�*( ^!'. a��]�*4 �'E ��/BI�u�7rI]�G�'��u�'W]BU�'��u�&֦�B�B::��B�"BҪB`8��]+z �!� �9���;��]+� �!'� ]$� �!� �9��ۥ ���,>�\� �����B �:%B �::A���-�$'� D�]���a]�������r�1G��]� � �!(��;�-��9��] E �!����!J�]���r�\����������\�/!�*�(� ����.]� 0!�!.!��-���� �-F]� H!�*F!] N!�!E ]="Z!�(�(�('�''m(K ]+h!�''�!]d$p!�(�W'|!]+z!�!'�!]�$�!(�W'�!M���B�B::'��:�/�!��Q'�!M��B�"BҪB�$"�P��]�*�!�'E ��E S���B�B�Q�!]�*�!B"�!�S'��]��]���B"ڥ���B�"B��B�]����E� ��E�ug'� ��E�up!�u�!�u�'Z!V����Q'*"�9��*!Y����Q'3"\���up&E$&"E]BC"gE� �\�Q�M"gg�9�����E ��Q'r"]$f"�!E _��:�:�E ��Q'�"�9�'�!V��9��'B�!Y��]$�"�!E \Q/�"�!�9���;-9ݱ�b��E e��E�u�$1�r�!�u�&E�'r�]"B�"�lqh��]�$�"('�"k�]�dB�"���� ���hZ&E ��� �-� ]O'�"�"�(�Tb��9��]d$#�(��]�*#�!#��;���u�&En��E ��]�$,#('1#q�]¿B72�E]��?2�E]�G2|���9���;�-�c�$"Ea9�.E w��'Bk1z�]"Bq2aw1}�]"�m�� *�m(�* &�����0 �`� � ��':	��O`eŅT��UTB׃ O�`�UL Q��Cg	 ,��Փ �S���4�g	,���]="�#�*�(�('�\!]s#�#g(�(��Ě��u"�1"E���E ����&B?� ��;9�;�E]��B�	A9�;�E;'�A�3'$1�'$�1�����]$$$�!)$��q9�;'�2�@��� �9A�\��CB�A]B�KB��rK����Ҩ"E]B_BeA�]rBkBvtA��xv1��]$z$�!�$�����]r���B|$"�A|�q��t6l'�l']8%�$�(&l']8%�$�(&�#�Q'�$����uv'�A�����Q'�$����u|'ܧ@;�r�]B���B|�A����|Q&E ;�&E ]�*�$|!E $E � ]="�$�*�*�(;��K ��Q'%����u�'Q�9�(%��Q&E $E ]�!g(�*��]���1R�;]R�;R����9���;�-�E�u�&E$"E]�g��Y� ]�*�]��K����@kPbb/bAb\b\R`�Rʎ�� :�Ш�� � �-�P]="�%�%�(�(x  �`�(�%��� 9� �` �`�%/�`M ���D V�`O``P	�# �� TRL� �0�H��9 r�'�ɔ3��I� ��� � �-�P]="�%�*�%�(;���%���%��� �1	��┎�� :��x X9�'��]RBbRR�]RBbgx]��#b^x�rUgRx]B5bp�]RB=bgR�Q�;�'�%3�'r��P+�'r�Q\��7%�%��9����Q��1�_%�%X� 9��s� 9�ߦB!B �:%B �::B�"BҫB\b��b�������\�/�&�*�(� �����`\�/�&�!�&��-���� �-�`\�/�&�*�&] �&�!�9����&\Q/�&�!�� 9�ߥ;-њ�9�;�-]���b����� �I!�]<r�'��9���]<!$'�!')�(9��|]<3r|'��9���U]<!B'U!')�(9��^]<Qr^'��9���]<!`'�!')�(9�����y]�<srX*���B!p]<!�'p!*)�(9��g]<�rg*��9���[]<!�'[!*)�(9��a]<�ra*��9���m]<!�'m!*)�(9���]<�r�'��9����;-ݦB]"���rB"�\rQ��rB!B�"B��B�]r��r���$��+]�!�'�*�� 9��]�*(�!(]� (�!(������I]B!�UI�&I�������;'7(��9����'?(��]��Ia�ڔ�U� 9��]$T(U!I!]�!I!�)]�!b(�*�'"m]��m�˥�����B!�}g�B ;\�(��qB%�'��e��qB%������B9�/򞙀��,B;��'�(9�'�(���t����7��B�"B�gZw(	R������(��,*'2'�(�������,:�(�������,�(�������,$)'�(����%}'������,zZ')�ԙ�wZ')�Ι��Ζ�;�n'� ����,�������,�����B��j�B;�r@����B �1���B�-B%j�0�*'"� 6���a�� �`� �� � ��/��O�`�T�D1�t�'�TX�`�DB#�t� '� S�N�!	l�����D� ��B!�m�B 9�B��B�"B�mZ�) �`�(�) �`�)/�O`e��$N� �S�Y��a8�@��*B:N-pY��2��p���BR0*B9���M� v������ v� �/���ȀE�%�X� 	R�RT�N�!ՃE�'	� ��O��Hɔ3�)���'B ����$ ����t�* �`�(** �`(*'��@�.*'Ӫ���* �`�(:* �`�*/�X�E�X(X 	�!RTN�� ׉�3`�`�T��@g��ϐ��4S	�S�gH��f�R�R]s2u�l�R�U]s2�`�R�X]s2��*�R�[]s2���R�^�a�]s#�.�)R(d�]s#�.$)R(g�]s#�.B)R(j�]s#�.�)R(m�]s#�.�)R(p�]s#�.W)R(s�]s#�.�)R(v�]s#�.9)R(y�]s#�.�)R(|�]s#�.u)R(�]s#/������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������     �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �	� ]ՠ4��C`X�	8��6A�tR]N��D�S ��F� �  �  �  � 	�( P]�c��D�`1EՃ	���Ag�RA]�N�T��@S� k  �  �  �  �	t ]ՠ4��C`X�	8��6A�tR]N��D�S ��F� �  �  �  � �� NL� �3�N�A`�1��TBRT`QX� ;�Dg��SRRQ݁��CA�4R`                      � (�p�o� &�n1�j�2�3�y�4&1�/67&5li���c3rDD��&%(/�ȯc5�$�/�k��n5�*�k��wr�k�s��2�/�5�7a.4/�4�3�n� �7!.5:&3�/57"5cc���5h/�4� ��!1� � �$�n%&f3�/5&5a.4�/2�/7"4@/ ��H$�!��!��k��d�֫    @ ^�h U@����c�X�$�(b� �@a��&�+%b&5bh���1�������5�/�5��n4/�4����4� ���3������ �t:�@H�1:�����:`"H��:d���`"����(:�(�2�(��3�b������֮݀�_)� �+�j^t)+�J� �!�+,&&/&%bib.�]b�%�(�J� �\t)�������� .:$f%&f���sx��%%���.��-��E��"��0� 	4�d����/�9��kilע�4��c�:�JccY��J74"P(��@�a4����&k �4�J����פ45&ccYks��i�8!.54&k��� �        ��1�/�5���/��+ $���k�5 @� �!��t)�J� �*��?��d        ��B�¨�Ӄ�� ����D��D��D ���b ���n��&����o��f�/��&�� ��b����&��0��&��3��@!�惃4��@��o��F���/��"J������݇�D �慢�/���� .��X���ƪ����V�������ݠ��������O�O���8�}                                                                                                                                                                                                                                                                                                                                                                                                ����P& � ]' �(O(���p9����dQ&. d;�-&�.� ��]�!6 �'�'B;��B"�������]��Ka�����ש��mڎ ;�&x \�-d (=(&j �:��:��:-� � :�1�^e%����m�V$"�|9�� ]�*� |!� ]�!� |!�(�B]"���B"�B 9�� �9�_9��B�-B�$� ]8%� �(�� "��̥  �\ *� �(\�+� g(j(m(p(�]�r�����!�����&!�.B��!�M!"pb�$�'U9���&!������6B:]B)�:�9�&:!]$8!U!'�'�E��E!�B\���Bŀ��]�$R!(�Q&Y!��]rs2ag���B]"s2km�����p�Y&�!��%�rB�u?"B� &�!��%B"���BR&�!��%�r�j��W&�!�����Y&�!\H.�!�(�!]�!�!�(]s#�!g(�*BҦ"�]Or�B"c��qB�&T+��,� ��2�""B\`������������¡��\�H�������\�H�"��� �]��"a�P�}�p9����"��Q&�!��Q&'"��q��t&x"� 2 �'l'l'�*? �*Y,x,l'l'E �,�.f/�/l'l'P!l'�!l'�"S#}#�#M$Y$l'l'W%_%\`-x"�(� ~ �'�(k*
+? 
+Y,x,�,E E �,�.y/�/	  E b!b!�!�"S#E E E �$%G%E E E \`-�"�(����;-���]"B�"�r�0&�!�&x" �`�(�" �` #'� %�8N X��5X'($@�]�"
#g(j(�) �`�(# �`P ''�@��uX&D1��,#�B,1��&0#����B>1��>#����XQ&�#��Q&c#�B!B ::X&[#:�B�!B�"BҪBM]2dBi2���&ru]2Bs2�&�]"�B{2��r�!�u�&�]2��2��1�9��#����"��Q&�# X&�#� �ݚE �^Q&�#]$�#a!�#a���"��Q�#��Q&�#�� &���� 6��':	���9 �T`N`�i)]��"�2g�j�� ���� 6�K�9y��y��&$\`-$�(��Q�+��Q�%��QS&��Qm&�����p� �9?�]�RAB?�L�BX�@�WX$�:�.R~a�r��/$]G+^$�'y�]O'h$y()��y�B�A�py�Tb��9�_&�$�:�R�\B`҉B���r��X$y�B�]B���B�&r�Ay�|$]+�$�'&�$|$y�$\H.�$y(|$]�%�$�'y��B��y��$y�M�]���B���y���y�y�y � �$%%\`-�$�(��Xy�\�+�&B]R��R�%���y]��R-��]��R��|A�9��&B}]R�-R����9��\�/8%�!�(��-�\���ER������ �9W�\��YR�WQ����� ���o�\��qR��o]RwR��y����9;9g;Xy�9�&�%�9�]����R��]���RE���9���9�]���R�y���;-ݨ9���9���Q���y���a��]r-��R�rڏP����������u&��]R��R��]��R�R�|�W6&��6&� 9y��]-+&R(&]�%&�'�W&&����p:�.)&��-�r�P��&6&]�!4&<)�+� ����F`]�%H&F&��9y��r/A�$^&]�!^&�(�-� ����9Eb����x&]�!�+�(]�!�+�(����.B�a��t�&��B�a��t�&�&���&��B�a��t�&��&B��`�¹a��t�&��&B��`���u��a�u�&��`����t�&��&B��`����t&�&њ]�!�&a(�+]�!�&�(��&"_q	�(�-��	�(�-�]�="r����롌	�-	%"m��m(�� ;��� ;�]�*$'U!,'U� 9�ߦ��p�WB�]�*:'B"P'��qB%U&H�p��]� P'B"�'��-��t/'���*]��er9�	�"	�m( �`�(v' �`�''	�΃� �NQ�E�"8�)�]�"�'g(j(�)�� v��� 6�P�;�l'3�&�l�pB�B::&��q:�l'B�-B�$�';�}�]r���r�&rE� ���u�&�q�9�6�'ܚ��Q&�'�9���&�'���Q&�'�9����p���p;-&E ��Q(��Q&R(]$(�!$(]d$ (�(�WN(���]�*.(�!8(�9����"�9���B(ۚ]�*H(�!&E ښE ���\�.B_]��]��K�ug&��g9�&�(]�*r(^!|(]�!z(�(K ]�*�([!&�(]�!�(�(K g� 9���gQ�(�[Q&�(g9���g[�}�]�^����]�^���r]�dB�����q�u�&?�r? �;�? ]�*�(a!�(�^Q&�(]�*�(^!&�(a��]�*�(�'E �gQ&c)]$)p!c)]�!)�($'g(\Q/)p!p� 9��]d$")�(���W&,)�����Q&:)�:)� ;��[Q&O)g9��O]��O�g��ug&[�g�9�]��K�r��u�&�]�Bo���\�Q�w��]���]�������K�ug&�]��������9�&�)]�!�)�)\Q/�)g!g� 9��p;9�;&�K���K ��Q&#*]+�)�!#*]�!�)�)\�/�)�!�(��-�\����������� �9��\������������ ����\�����]�����9����u�&2�m9;Z&:*]�!8*�()�� 9��]+F*m!N*�� 9���9�����]�!^*�!�*�9����;�-���r*����]s#z*g(�*B��B��B�$�*B�Y�*B�Y�* �`�(�* �`�*'��l&"�)]��"��g�j�� ���� 6�K� �͖r�Қ�]$�*y!�*y��]$�*|!�*|��]+�*j!�*j��]+�*X!�*X����*]$�*�!&l']$ +�!+����E �yQ�+�|Q�+�jQ&+����uj&/�j9��B/̰���u[&8�ؚ��RQ&A+����uXM��u�&P�ޚ���&�E]B[�RE�u���"v���!&q+�� !�B X�9����qX�9��u�&��X�9��X�9	��}�rB� ���|Q&�+��q����|]�*�+�'�+��7�]������&������|��Q&�+͚��&�E\Q���y]���|]�����$�E�u�%�횜�9�&� ���9�&�	������Y&E �9�;�-Ѭ9��B��9�ߧ9�;�-�E��9��2�᚜9;Z;,�����Y&E �9�]���I��S]��S����;�-�E]B_�UE����.EU�9�]��s����%*/K ]$~,U!E U� 9��]�!�,�)]8%�,�(K ]�!�,�(K ]�*�,�'&�,�^Q&�,]�*�,a!&�,���^Q&E ]+�,s!E ]�*�,�'E &E s� 9�_9��s� 9�_��]�!�,s!�*K �B!B ::X&�,:�B�B�"BҪB��B��&�-B-���]$-p!-���p�]r�%Ҡ5Ѡ9�&5-�����]r�;ҦDі�x�1��]$J-�!Z-�9�&�Zі�x�1����6Blq�&r�]�Bi�guџu�&u�g�]rB{�y&�]�B��|�����y1����6Blq�ug&����$&E \Q/�-g!g� 9��p;9�;&���������&r�����yQ�-�|Q&�-����up&������Q&�-���u�&��$'"g��u�&������Q&�-���u�&�9���&T+:���u�&E�9�&E ]�!$.*��}�\r��5�g�j�m�p��Z?.�&��]�G�����9����9��9;9g;�Tb��q����\�/l.�*�*��-�\���y���\�����\r������p����;1;Z�.;1g[&�.\�/�.�'�'��-��t�.������#��Q�.�&�.]d$�.�(���l']�*�.�'E  ���u���u�&E��9��p�;�#��]+�.�!&/]+/j!E ]+
/j!&J/&���u�&E�9��-�]��%����9��-�]�Or5���9����1���T+9������#j� 9����Q&\/j� 9��j)9����E ]$l/�!l'\Q/t/�!,��E�u�n�ug��up��uy��u|��u���u���u���u�&E̚�E �&�/]�$�/(�Q�/]d$�/�(�Q&l']$�/�!l'��/��Q�/Y���YZE ]d$�/�(�Q&E ]$�/�!E �� 9���   /    ��!E2M%*��:ѦB\" �����\ @ `�(        �-� E M A  ��������-�܂ O�\��SO���,\�/-    �     � �@FE` Ml m ::o.��:q:�p9y�@ `  ��' f     � �ЀE`MlA  �Ȃȃ��5B��� <� � �\�-\���u%� ����� �����R����� �����  !  � 8E� M� � �R	�p�:q>*   @ `��M�\r �  (� �ЀE�M�A  �Ȃȃ��5B&�� <%!!\�M\���,!���-݃����}������ g!    E E�>MIJg��Q%Y-�  9;�j��1;Z  C!     �e�E>!MI!A  ����������\�/�!�!�!��e!�!   DKE�M��U�-U1���/.�   @::Qo.\H.�-  �!    o0)� �рE�M�A �Ȃȃ�\��-����������,\�.�!�!�����$�!�����,�Bֆ��LY�#�!�!!"   �DKE�M""	�r]����r]���r"� p�!     �� E�!M"A  ������ ��Y2""�   E� HE?"MJ"K":*:%:%o�ঋ, -\.  @  bc) D     �Z-o.����BE&� H` h ��  �� 8 ��f"� fҀE?M"JA  �ȂȃȄ��"� ��]��"�\"���"n"_"_"_"_"_� �B܌ �B܌ �B� �B� &�\"� &��/*��A���ŠT`QUSA	�S�@����}� � ]�!}"�"��}� � ]�!}"�"'#   uqE�M"	2
2/���q'+��MQT�Ճ     ��]b� #     �%�0E�"M	#A  �������������I# �`#n#� � ���BX 6�2e�1 �` �` �`#j#� � �%':���)�'���'�,�)�� 0��� Eu#M�#�#"�A�/]"c��U(     @
�  � p z 0(   � p@    P  � �#� �ӀEuM2�A0 �Ȃȃ� ����<���#�-֋0�Tb��%�#��R��0��,Z�#\`-�#�#���-� 6��2�A �` �`\`-�#�#���-�]2OrB�2��<�#'�Y��=H'�)�B @ � HE$M$$%$nR� 0 UU!  � �=A�   @   � @ԀEMB$A@ �ȃ���Xa$��a$@�@@$�$   	`4 E�fMBqBr�D�$�B�@  @     @             k$     ���@Ef$Mq$���� 	�_�	����]�'�$�$�$����I����T+������"�B� @ 	L�CE�$M�$�$RR      @     P  ( � @            � �ԀE�MB�A@ �ȇ�	���T+���]O'%�$�$��L	��Tb��]O' %�$�$���B҂B)��B�Tb����1����$c%   � E�:MRERFnUp%�� @  @     ` �Y� ]� P  ?%     �a�PE:%ME%��]$t%U!}%U	�%�Q�� �-�P]O'�%�%N%%�%�aPa%�%   �U�E2�MR�R��U�% ` `  `
�   �.�r�uV�`   �%     ���PE�%M�%A  ������� �-�P]O'�%�%�%� ���5�������P�-      �>b `��D�A�5;ցg8`Ai8�d-0&��A�M�aD`>-*&;�%5;v�%�;b`  @  
   @�          �`!G&Ib��Wa�`Q&�]bZ`\&���d`f&�:5�n`p&�3-�x`z&       �R �EB�Mb� `                ��R��]�#�*    �& �b�`���`E�&M�&A ����ȃȂ��Ub�h P�ҫUb��a !��&E'C � ���ׁ�WA 	 B  ����Mtqt-r�`p pЁ�u�&�&      ECp � `          OMp� 8E/'M,'      
� UP]<%B+U%'-�,  ( p( ��Hp�H�pE/'M,'A ���������J5rfp���5m'A  ��=bJp��yGHEr�Cp �����q�E�Ap	  B  Ё���M�G��G-�' �'  (�����R�r� p � @E�'C  '            �`  �` ��0<-ѦB]b����Bb�]�Q2��BaB�bB��B�]��R�����$��/]�%�+�.�� �*9�&�	�������EE"M�� �a+9��@@ p9�ߧ9�;�-�E��  ( ��\9;Z;,�����Y&E �9�]���I��S]��S����;�-�E]B_�UE����.EU�9�]��s����%*/K ]$~,U!E U       @     `     P     p   � @   � P   � `�    @@  � @   � P�    `@  � `�  @ p�    @`  � @�  @ P`  @ `�  � `   @ p`  � p�  � p  ` @    P   � P�  � P0  @ `P  � `�  0 p@  P p�    @   @`  h @�   PH  P P�  @ `h 	 � @	( 	 � p
� 
 � p � ��, N  ( : %! g �-- � p�  � �E& � p, \ ��/ y ��) 4 @*" ; ��/ r  :( � P�.N �R X��T ��  �� � ��  ��   Pp  � p   � `   � `�  @ @�  � p�  X P   ` Ph  � P�    PH  � P�  � P   8 P�  ( PE�d `�  ��  � @    p�  @ P�  � @�  � @   � P�    P�  � PP    ``  � `�  p `@    p�  � `�  � @�  ( @0  8 @x  � @�  � @�    `�   `    `�  ( `0  8 `H  P `x   @   � P�  � P�  � P�  @ @� �  ��  � @  /��/��E(M(_ � E�A�  �ȱ����� �\UJ&E(]+a+E�*A  � )�ȁ�����U�J�l-XUJ&�U"QEb���"aE��A�  �Cȱ����� 	��UBJEb��aE��A�  �]ȱ����� 
��TbE�j�Y \ �g����]="s� ����;���py���;��+��+y�+�B�]����6��y�!%"���Ҧ!!y���]�-���%��\��ҷ���%�ۦ�B�B:*%y%��:�%���y]������B�"BҪB��y��*]�-���%�*\�����y��%�*�:%���-*/�:*�:�%b,�-B*\�H��%�*��:ѦB\" �����\H.(,�(0,� ::�B�-B�$,�B!B ::X%H,O::�:::*�B�-B�$;,]�!Z,�(]� */�!(���̦B!B ::o.��:q:�p9y���,]�%�,�'y��5B��y��-�,By:�*"����t�,y1�:�����t�,y::Q�,]-+�,y(%�,B�%B�\�����y��%��]�G�����t�,�y9�:���r����-�t:�R~��pB:*1-:���t-�,��M�\r ���r��:::*��1::�:��--:%%%-::X%-:*X%-�&��:%�o.::�B�%BE��"o�9�o.���p���g���Q%Y-�9�;�j��1;Zj-]�*h-�'%�-]$p-�'u-��q��r��gZJ-��%�%�ќ%r�Ѿ;%�-]$�-U!�-U1���/.� :*::Qo.\H.�-�(o.]�!o.0)]�!�-3)�;%��\Ҕ��Ҿ"\���ү%����j���Q%�-�9�;���1;Z.]+�-�'	.�;-%�	]�^	�r]����r]���r"��r��jZ�-� "::�:*ҥ:%o]��5�N\���=�"\��"�%���,B:*:%:%o�ঋ, -\. �\ *b.c)��:��H�Z-o.����B�"BҫBi��*/�B� ������ �` �`�./�RQ`R`�q'+�A��3T�`QR��TN(�),����CT� O&n�Y]�!�.�(�*�:�%�.�:��B ����ҋ� �` �`�./��q�'��M�#����TT�g8@���כ�5�.��-�]���∛�*// �`�(/� � �/���q'+��MQT�Ճg@����]b�%�ǀ���.�&:r-�p��"O��� �-J�]O'N/J/"���V/�%]/:4M�]r-�c�%�~]�8Rk��~��x/\H.v/�(&�&� ;���]�*�/�!�/]�!�/?)Y�#�/�'��]r-���&��1��%�/\H.�/�(�/%�/]�!�/�(]8%�/�(&K 9E�b9E�;�B�BK ���B���t��dQ%�/]�*�/�!&6 �9��$&"6� 9����Q�/��Q%�/�9��
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
 
  P
 
  P
 
  P
 
  P
 
  P
 
  P
" 
 * P
. 
 2 P
6               
8 
 : P
< 
 > P
@ 
 B P
D 
 F P
H 
 J P
L 
 P P
R 
 T P
V 
 X P
Z 
 \ P
^ 
 ` P
b 
 d P
f 
 h P
j 
 n P
p 
 r P
v 
 x P
z 
 | P
~ 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
 � P
� 
   `
 
  `
 
 
 `
 
  `
 
  `
 
  `
 
 " `
$ 
 & `
( 
 0 `
4 
 6 `
8 
 : `
< 
 @ `
B 
 D `
F 
 H `
J 
 L `
N 
 P `
R 
 T `
Z 
 \ `
^ 
 ` `
f 
 h `
l 
 v `
x 
 | `
� 
 � `
� 
 � `
� 
 � `
� 
 � `
� 
 � `
� 
 � `
�                 �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �
�  9�     �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �	� ]ՠ4��C`X�	8��6A�tR]N��D�S ��F� �  �  �  � 	�( P]�c��D�`1EՃ	���Ag�RA]�N�T��@S� k  �  �  �  �	t ]ՠ4��C`X�	8��6A�tR]N��D�S ��F� �  �  �  � �� NL� �3�N�A`�1��TBRT`QX� ;�Dg��SRRQ݁��CA�4R`     @     @     `     p     @     @�    P�  � P�  � P     `�    p�    @@  � @�  � @�    P@  @ P�  � P�    `@  � `�    p@  @ p@  @ p@  � p�  � p�    @   @ @`  � @�  � @�    P   @ P`  ` P�  � P�  � P�  � P�    `   @ ``  � `�  � `�    p     p     p@  ` p�  � p�  � p    @   0 @P  ` @p  � @�  � @�  � @�  � @
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p
� 
 � p     @   @   @   @   @  	 @
   @   @   @   @   @   @   @   @   @   @     @   ! @"  " @"  " @#  $ @$  % @&  & @'  ( @�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � p�  � X�  � X�  � X�  � P�  � P�  � P�  � X� �� P�  � P�  � P� � h � h! �# `% �  �                           �D@ 	� 8N P�� H� ��� H�� π� 8��5 ��� �E �� X�S ԄI � 5 Ճ XXT �V �L �S X� Ԅ� H��@ ��  �W  π� N�% N�� HN ( Մ� H�3 ��� X� �� H�S �� X�� W�� (�N ��W P�U P�  �` X B�� 8S�   �  �� �� H	 E Ճ X�C  ԄP E �� ��A � 8�P# ��� H�R1 C�� HA� `�  ���T ��  ���4 ��  ��TE ��  �� 8 ń  �� H ��  �� � 8�S ��� 8r h ̀M (�3 X�M CU �� H�� ��� 8�TB ̄B �f � HN �G X��@ ��� X�� �� �C ҃E (�� ȄL ��D A�N (Ɖ1 ��� H�S& ł` hP3 �D �3 ҁT �� ��  � A ԄP �� �� 8	C �� 8�K@ ��� H�P ̀M ��4 A�� S�$ ЄL �� �R �F" ΂V (�� ��	 X� ��� H�U 2�� 8� 3 I�� HN@ ��N N@ ԄL �D@ ��� X` �W 	�D �G �S  �� 8�S ��R E�4 �� 8�S A�� ��S �� X�� O�� H� ��� 	M Ʉ 8�� ��� X�N ȀS �  �A G� G�� ��4 �D (��T I�� 8�R@ � XMR �T �D �R ��A �� H�CB ȀI �� �� (�P! �� X�AA �� H�  � X� �� 8�E 	�� HP ��` h�N  Ʉ� 8TU U�B 8NS ЃN �5 �� �� 	�� � 8 X�	 XƠ1 ��� X�K@ ׄN (� �C ES �� 8��C �V �  �� 8ϔ X� H� �� 8�T T� X�# ��� 	 % Ԅ� HRE A�  X� �N (��@ �� H�T U�T (�� ȅR N�% ��D � ��S  G�� 8�� Ä� 8�` ��` �` ��� 8�` ��E (�D@ �� H�A ȄT �S@ ��� (	� Մ� HSE ��� XR% ��` �` ��` �� ��` 8��D ЃN B� B�� H�Z@ �� �@ � 8� � �E EQ 	�� X� �� HI�4 ȄT (N ��� ��C N�� �MB  �  �                           	� � ������     �*�� E�!M"� A D�"L�3�4���Y2""�  E� HE?"MJ"K"X  -*    ���(�b��         � D  (         @     `
�  -v
� � O*� OڀD"L�3A� �������$����Y�B��l�����\�����`���Tb����\����c������T����*�*�*   �L@ D2�L����Ť��ŠTP       @
���}� � ]  �* ���뀠D�*L�*�A�����������,2�� �Q � �D+L++  � 0# ��%�0E�"M	#A  ������  �        @     @   @ p  � ��:��D+L+A  ����������������m������������\�`ҁ�K]��b��0�?�3]��b��0�<�0]��b��-�E�-]��b��-�B�*]��b��-�?�']��b��-�<�$�Ѓ�Є�:�)��<���#��	�SD�+L�+�+��R��0��,Z�#\`-�#�#���-� 6 � �    �` �`\`-�#�#���*;�A;'� ��EE" �        `     `    !-  � �����D�+L�+A  ���ȂȃȄȅ ��I ƆK1�) f��]A�� ��	`L�S Ɔ`2�i̓��������������4K,� <!�Bj����,�����4�,� <!�$Bw����,�4B���<!���,���������,�4B���<!��$�,]'�,,�+�]�r��������� � �-��]�&�,�,, ,� �<!�Д�,�B������ ��\����������$B��'�����!݋ ���@4!<!݋���!����Ѕ �\������'�'�� `�  0 p@  P p�    @   @`  h @�   PH  P P�  @ `h 	 � @	( 	 � p�-   �� D�bL�m�n�N  ( :   g �-- � p�    g-     ����Db-Lm-A  ����� �`v-�-� � �X�(��� SR���Is'+ ϰ�L5 OVRX�L0Z�R.�@�. 	 �TD�L������,   (�p� `       @�   �- �  @     @     @     @	  
   @     @     @     @   ���D�-L�-A  ���������	����>.���T�����T+���UQ&�-s.    E D�JL�U�V �`  � `�   @ `    p�  � `O.     �q��DJ.LU.A  �����\ *�.a.�R���q.q����   `  O  �D�.L�.�.0  8 `H  P `x   @   � P � �   �  � P�  @ @  �  ��  � @     @     `   � `�  h `   �/ �������D�.L�.A  ���Ȃ��Tb�����&/ �`�.�.A� �`	�LO �`�����]�Or3����蒍,� <Ғ�� ��4<-���,�B>�����| � �SDS/L^/_/ _\� �    � ];"s� ����;���p X �z/� z߀DSL�^��A ���\�/z/�/d/�/   O�5 D��L���y���]�-���%��\�@ 	 � @�%�� ��/     ����D�/L�/A  ����������4�/�����-�����4B����]^ �/�/�/�  ��  ]� �/ �� @     P     P     `     `     `   � J�  � P�  � P�  � `�    p� �� @�    `     p     p� �� @�  � `�  ��@�� ��@�    @   � @�  @ @@  @ @�  � @�  ��@�� ��@�� ��@��   p@    p�  � p�@IPgKP�KPkKP�KPk�  � p�  � p�  � p�  �@O�@�PO�P�`O�`�  @H p k�           � p0  0 @@  @ @@  @ `
  0 @0  � P�  ��Q�  � P�@IPgKP�KPkKP�KPk@    P   � @�  � @     @�  � @�  � @�  � @�  � @�  � p��0� P�    `   @ @@  @ @`  ��H@    @   � p     @   � @�    p   � @  � @�  � @�  � @�  � @� 
 � @
� 
 � @
� 
 � @�  � @     @    @   @ P@  @ P@  � ``  � p�    P@  ` P�    P@  � P�  ` P   @ `   @ P`  � P�  p Pp  � P�  � P�  � P�  @ ``  � P   ` `�    `@  � `�  @ ``  � `�  � ``  ` `�  � `�  � `�  � `     p�  � `�  � `�  @ p0  @ P     p�    P     P�  � p�  � p�  � p� � p�  � p�  � p�  � @�  � @   @p  p `�    @   � K@  � K �� @d `� @p  � K�   @0  � K�    `+ � `   � P�    `   � PP  P @  @ @@   Wp  � `  p @   @�   @`  � `  ` p�   `  � @�  � @�   W�  � @�  � @�  � @�    @   � @   @ P     P    P   � P�    p@  P P   0 P   0 P0  � `�  � P�  @ `@  @ `   � P�  @ `�  � P�  � P�  � @�  � P�  � P�  � P�  � P�  �pF�p`�pF
�  � P�  � P�    @     @�  � @     `    `  0 `     `	� 	 � @@ 	 � @	� 	 � @0  ��H   P `P  @ `@  @ `p  p `p  ` ``  � `����x   p `p  � `�  � `p    @  � `    @(  0 @8  @ @H  P @X  � p� � Q� � Q� � Q� � Q� 
@� @P   p  p @   ` @� �� I� ��b�   @   ( @0  8 @@  H @P  X @`  � `�  � `@  @ p0 
 � @`  !�w!�p!�w!�pPW	�  P_
�  � @P  P @P 
  P
  P @�  � @� 
  P
  � p!�p!�w!�p!�w	� 
 � @�  � p  � p�  � p�   @�  � p�    @     @�   @�  � p�  � p�  � p�  � p�  � p
� 
 � @�  � p�  � p�  � p�  � p   @  � p     @�   @   @  � p   @�  � p�    @(  0 @8  @ @H  P @X    p�   @(  0 @8  @ @H  P @X    p�   @   0 @8  @ @H  P @X    p�   @   ( @8  @ @H  P @X    p�   @   ( @0  @ @H  P @X    p�   @   ( @0  8 @H  P @X    p�   @   ( @0  8 @@  P @X    p�   @   ( @0  8 @@  H @X    p�   @   ( @0  8 @@  H @P    p     pA@K�F���dP�@�?�M���� ��F����������&��?���
� 	 � @            �   � @                                        O�A��L0L� �CDD L�1 N2 E��  N � �$� 3XL`!�� p                                  `p    @            p�         @ `�               @             `  � `�  � `                  �                                                                                                                                             �                                                                                                                p     � @     P@           ` p�                    @         �  � p�                               �          @              � @�           ` @                                         � @                                                � @                                  P         �                                                                   @      �    @                                                                                                                                                                                                                                                                                                                                                                                                                                                       ( @                                                                                                                                                                                                                                                                                                                       `     P�         � `�    `�  @ @P  p `     � `              `         �  @ `�  � ``            p  P pP            �  ` @       `                                         � @�    p@  � p     � P�   `@  P `     p p�   @                                                                                                                                                                           �               �                � `                                              �0    ��           ��  � p�           �     �       �                                                                                               � p       �                                                                                                                                                                      	 � P	� 	 � P	� 	 � P	� 	 � P	 	  `	  	 ( `	4 	 D `	P 	 X `	h          	 p `	x 	 � `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	 	  p	0 	 8 p	L 	 X p	` 	 l p	x                                          	� 	 � p	� 	 � p	� 	 � p	� 	 � p	� 	 � p	� 	 � p	� 
   @
                                                                                                                                                               
 
  @
( 
 * @
. 
 0 @
2 
 4 @
6 
 8 @
: 
 < @
@ 
 B @
D 
 F @
J 
 L @
N 
 P @
T 
 V @
\ 
 ^ @
` 
 b @
d 
 h @
j 
 l @
n 
 r @
t 
 v @
x 
 z @
| 
 ~ @
� 
 � @                                                                                                             �     �     �     �     �     �     �     �                                                                                                                                                                  �                                                �  � p   � p     �`  � P�  � `@   ` @                                � @�    @�    @   � @     @     @     `     @�    P�    `�    p�    @@  � @�    P@  � P   @ `   � P�    @   @ @`  � @�  � @@  � `�    p   @ p`  � p�  � p     @   0 @@    @�    `   @ @�    P                                         �  @ `                        �  ` @�  � @�
  `P  p   h `   ` @� 
 � `
� 
 � `
� 
 � `
� 
 � `
� 
 � `             	 � @	� 	 � @	� 	 � @	� 	 � @	� 	 � @	� 	 � @    	 � @	� 	 � @    	 � @	� 	 � @             	   P	 	  P                               	  P    	  P	          	  P    	  P                                                                   	   P         	$ 	 ( P         	,      	0 	 4 P	8          	 < P         	@                                                            	D          	 H P	L          	 P P	T 	 X P	\ 	 ` P	d 	 h P	l 	 p P         	t      	x 	 | P	� 	 � P    	 � P    	 � P	� 	 � P	�               	� 	 � P	� 	 � P	� 	 � P	� 	 � P	�                                                                                              @     `   � @   � P�    @�    P   @ `   � p`  � @�    P@  ` P�  � P�    ``  � `�  � `   @ p`  � p�    @p  � @�  � @�   P@  P P`  p P�  � P�  � P�  � P�  � P    `   0 ``  p `�  � `�  � `   @ p`  � p�   @   ( @@  H @P  h @p  x @�  � @�  � @�  � @�  � @�  � @�  � @    P   8 P@  H P`  p P�  � P�  � P�  � P   `  8 `@  H `�  � `�  � `    p`  � p�  � p�  � p�  � p	  	  @	 	 d @	t 	 | @	� 	 � @	� 	 � @	� 	 � @	� 	 � @	� 	 � @	�                                                      � P@    `   � @`    P�    p�  � p   � P`    �     `   ` P�  � p   � P@
    `�    @�  � p    P 	    @   � P   ` P�  @ p   � P�    ��  ` P�    `   � P   � P@
    @�  � @`  � P�    `@
    `   � P   ` P�    P�    @�  � p   � �   ` P�  � P     @�  � P   � @�    ��  @ p�  @ @�  � @�  � p�	  � P   @ P`  � @�  � P`  @ ��    @@  � @�    ``  @ `�  @ p�  � p@  � p   � p`  ` `�  @ p�  @ ��    @`  @ ``  � P�  � ��    @`  � P`  � p�  @ @�    @�
  � @�    p�  � P   � p�  @ p�  @ @`  � P`  @ p 	    ��  ` P�    p   @ P�  P @�
  � @�  ` �   @ p`  � P�  � P�  � P   � P     `�    �     �`  @ P�  � p�  � p�	  @ p�
  @ p�    p 	    ��    p   @ P`  P @   � P�
  � @�  � P�  � `�  � ��  � P`
  � @�  ` P�  � �     �    @�  ` P�  � `�  p @�  � p�  � �`  � `   ` P@  @ p�  � P�  � P@  � p�    �   @ p�  � p   � p     �`  � P�  � `@  � �   � P@  � P   ` P�  � P�  @ p�  ` P�  � ��  � P�
  ` P�  � P`
  � P�  ` P�  @ p�  � P�
  ` P�
  @ p�
  ` P�
  ` P�  � p@
  � P@  ` P@
  � P`  � P@  � P�  � P�  @ ��  � ��  � P�  � �@  � ��    p�  � P�  � �`  � �   ` P@  @ @�  � P�  � �`  � P@
  � P�  ` P@
  � P�
  @ p   ` p�  ` @�  � @�
  ` P�  � P�  @ p@  @ p�  � P�  � p�  � P�  � P@  ` P@  � �`  � P@  � p@  � P@    p`
  � p�  � P�  � PP  � P�  � P@
    `�  ` �`    `�    `�  � P@  � �`  � P�  � ��  ` �`
  ` P�  � P�  @ �   � P�  � P�
  � P�
  � P�
  � P`  � ��  � P�	  ` P�
  @ p�
  @ p�  � p   ` P�  � P@	    �   � P�  � P�    ��  ` P`
  � P�  � ��  � `�  � P   � @`
  � P�  � `�
  � P�
    `�  @ @@  � Pp  � P�  � �@  � @`  � P�
  � P�  � P�  p @p  � P�
  � Pp  � ��  � @�
  @ p�  � p�  � P@
  @ p�  � �@  � P`  @ p�  � ��    `�    `@  @ ``  � P�  � ��  � P�    `   @ `@  � p`  � ��  � PP  � P   � P�  � @   � p�    `�  ` P@    `�  � P�  @ p@
  � P�  0 � 
  � ��  � �     P@  P @�    P   � @   � p�  � P�  ` P 	  � P�
  ` P�  � P 	  � P   @ PP    `   � @�    p   � P`  � @     ��  � P�    `�  � p     ��  � @�    p`  � ��  � P�  � @�    ��  � P@  � @ 	  � P@  � @�  � p     ��  @ p�  ` P�    P     ��  � P�    ��    `@    `�  @ p�  � P�  � �@  @ p�  � P�    `�  ` P�    �@  � p�  � P   ` P�  @ `   @ ��  � P@    ``  � p�  @ p�  � ��    `�  � P`  � P   � P@  � �`  � P@    `�  � P@    `�  ` �   � P�  � p@  @ `�    ``  � ��  ` P�  @ p�  � P�    `   � �   @ ``  � P�  � p   @ p�    ��  � �	� 	 � @             	   P	 	  P              @     `     `     @     @     @     P     @     @     @     @     P     @     @   � P   � @�    @     @     P     P     p     @     @   �j���j     P     @     @     @     P     @                                                                                                                                                                                                �� �ɴ&˼&�!.��s�.��r��r��b�F����s��r��s(����dǁ<�|ǟJ�̄.��/��0��1��� ������堛� ����֐�נ� @E � �   ����� � � �����                                  @ ���"H�����"�����B��t��"�����&��˃��6 ��/�����n��&��B��/�����b��˂��0� ��~�      T                                                                       @     @@             @@�� ���?�����i��ω������i����������i� ω�� ��҈� �ޢ��b��&��Ɉ��
ܺ&��������/๜�����������2�����ˑ��̄濊����d���� �������  8  0  (       � � �    @   ��&��� ������è�/���ҫ���h� ���������� 𗭢��h� �� � ��(�������JB���6��Cвd��6��Cϲd��6��LБ<��t �� ��É�� �    ���bЁl��2@������0��'��J��˝x���� @������h  �����     P     @     @     `     p     @     @�    P�  � P�  � P         �  � @   � P�  � P�  � @�    P@  @ P�  � P�    `@  � `         �  � @@  � P�  � P�  � p�    @   @ @`  � @�  � @�  � @                                                                                                                       @     P     @     @  
 � @
� 
 � @     P     P     p     p���J�
�� @� �� J
�    P     P     p�  � @�  � @�  � P�  � P�    p�T �8� ���#   �AA�A"�I2�2��;������� ��  � � �����  ~ (����  �#    �0���0A�#I�#A  ������=�0��\2���2�1��#�Ȁ�A��-\�.�#�#�B�2��9����&�b�l���Jj�����T���7�- Ww&63��9	�� A;$� ��⟁l��'��$��rF$��|� �� !�@ ����O� �  �  �  �  ��A���d �� �   �G �S  �� 8�S ��R E�4 �� 8�S A�� ��S �� X�� O�� H� ��� 	M Ʉ 8�� ��� X�N ȀS �  � ����b��&��&��ð�/�������⪋j��&��ë�b

�
�諲(��D���Ń�� �   
 #���q � �(/��(���H/��"��Ȳ���&� ��l���ׁl��?��D���H/&���ŉ����)��?� @ ��`�T � ЃN �5 �� �� 	�� � 8 X�	 X �܊&ږ&ň& � ��.���@��

�
�� ������*       �������b��b��b� `� 0�� � ��.���@����.�  ��|������ ��� ���&�� ���& � ��.��@�➘o@�� ���&�?����   ���o ��` �`8&� 8�` ��E (AN2 A��IR�R��TD&�S@ ��� (	� Մ� HSE ��� XR%  ��%    �` �� ��` 8     `     `     P`  @ `�  @ `h 	 � @
�   E& � ��& � p�, N  ( : %! g �-- � p�  � �y(  0�! � �4$ *  ;*  ��/ \ ��/ r  :( � P�.I�%A�%Y $Y  ]�']�'X� X�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
� 
 � P     �   ` @@   @@  � p	� 	 ( P	t  � N  � @
� 
 � p                                                                                                @ @�  @ @�  � `�  � @p    `�  ` p�  8 @�   P  ` Px  � P�  � P�  0 `@  ` `h  � `�    p(  8 p@  � p�  � p� 	  @	$ 	 < @	@ 	 ` @	t 	 � @	� 	 � @	� 	 � @	� 	 � @	� 	 � @	  	  P	 	 $ P	, 	 D P	L 	 P P	l 	 x P	� 	 � P	� 	 � P	� 	  `	  	 8 `	H 	 T `	h 	 t `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	� 	 � `	 	  p	 	 , p	8 	 D p	` 	 p p	x 	 � p	� 	 � p	� 	 � p	� 
   @
 
  @
 
 & @
: 
 @ @
D 
 P @
d 
 j @
l 
 n @
r 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 � @
� 
 
 P
 
 & P
: 
 N P
b 
 v P
� 
 � P
� 
 � P                                                  `     P�         � `�    `�  @ @P  p `     � `              `         �  @ `�  � ``            p  P pP            �  ` @       `                                         � @�    p@  � p     � P�   `@  P `     p p�   @                                                                                                                                                                           �               �                � `                                              �0    ��           ��  � p�           �     �       �                                                                                               � p       �                                                                                                                                                                     @ p       @       @�  � @@    p`  � `@  � `�  � @@  � ``  ` pp  � `0  � `�  � @  � @�  � `�                      P     P     @     P@    @              @                       @     @                                     @                                            @     @@  @ @@    @     @     @@    @@           @                                                                                        @     @@             @@    @       @                       @             	   @	 	   @                           
                       @       @                              @     @�    @     @                                                                                            X� �� N     P   � @@    P  � � @]�cV�`C	V!D(TN�"�Xg�DN� �D�u�R5R�͐z�F.��o�<��t�����(�����r��~�� q    !ϥ���?���D����&��!�ʀ���(?ސ���É(��Φ����&��&�� ���9  �ͣ��I� �
����"Ͱj ���&杯x�?������ ���2@������0��'��J� ����������������                                                                                                                                                                                                �� v      ����H����   � ��      ��� � ���BD `       	   �         �     �Ѐ ���8 ��#��� P��I� y4�� ������������0F	 q�*�=���c  ��+��/.
 A�5? ��a\ �� T �8� ���� ����K���������������� ��   !�L��� {�~ (����!.��/�����޵�ҷ�cH������v� (��� ��B���� �����H��k�(������Ť)D��H/&��ˋ������&�b�l���Jj�����T���7�- Ww&63��9�nӇj ��i��̪�̪̱�����?��CH�(� �����̏�!��"�`&��X��j��},���̀������;�/�ӢD�� �����	��}�
�̳����D.Ҥ, �    ���l��&�����rD�₁��˒�'��&��& �&�|���&����d����'� �   �� �~�{ �zіz��6fy��c00b�:f�0�x�����/u�/n�/r�/c�/������ �/� �/�9�:b(� �:dw ����������ɼ��0H.@��n�)˩l0.����:F.:D.9�*�" ����'w�/�&0':(/!��w�������/v���������3"[�(��"��h��u�����0uI��/������� ��/�u�t��s����r��bF��⩕�'�0ē ��$����:&13f2b���"���x)�����f����� ���������������� 	�q����p��q���:��!N6�n�j�����:&����gp��;)�a��"9V�9��@.o/������@O�9����9�c��o���nIH.����v����%�b&�h��sV��s��m2�t�y�!.li�Ȩ��8t������
�

�r��"H.��&��!8���y����H�����J2����L��Ɉ �
��� ��2zyw�NziOkiN� � �6d3G$0 Ə/v��j�i8�`o�����H/H$.����2 H��2HHb&��8D.8�"
�k� ��H����H�HBbhC�D�Fpk��H$.����H�HFbG�h
7�Jk�B��<�
�b�b�k �t)@�/����t)C~ D.����k82F�8(/��"<�h
7�JB| �J&@�+�����?��:{ �@�/gھH����C~"Ih!>FF&p �`F�Fo�C�f����$����8��eb��kU�_CC4 d���/p����Bh !C�H���D��Cf�H�H��H�nf���тDDb�/�C�C�i�Ѩ�h�Ch0�CdCh0J
�J.
��    �C�                               � (�p�o�,&�n1�j�2�3�y�4&1�/67&5li���c3rDD��&%(/�ȯc5�$�/�k��n5�*�k��wr�k�s��2�/�5�7a.4/�4�3�n� �7!.5:&3�/57"5cc���5h/�4� ��!1� � �$�n%&f3�/5&5a.4�/2�/7"4@/ ��H$�!��!��k��d�֫    @ ^�h U@����c�X�$�(b� �@a��&�+%b&5bh���1�������5�/�5��n4/�4����4� ���3������ �t:�@H�1:�����:`"H��:d���`"����(:�(�2�(��3�b������֮݀�_)� �+�j^t)+�J� �!�+,&&/&%bib.�]b�%�(�J� �\t)�������� .:$f%&f���sx��%%���.��-��E��"��0� 	4�d����/�9��kilע�4��c�:�JccY��J74"P(��@�a4����&k �4�J����פ45&ccYks��i�8!.54&k�����        ��1�/�5���/��+ $���k�5 @� �!��t)�J� �*��?��ds���	&�js��n����^t)�s�x����_��_� P���H%�&n$d�y� .li����)%�/��"t��!.b���"H���n���*�j^"���s���	&���t��η�eb�! �����| ��&� �&�
&h�&�Á
���Je� �n�;�͸����I����p �H X�R(	�H��(��r�^&��@�"�����h
o��n@�/�@�dx	�L��4��.��N��C� 9m@/ԗ��	�w����!.��0����\��	�	�n&��(�Ȗ���|	���	�h�
-^b��h0�	tԼ�R�c� @ޛ �����f�IC�C N���fIhD�K�D��C�C�d���ѓ 0� ^@r���&�/�֮A���xO��Po�Uo� `�@���/�o��n�b9�n��&@�/��@��9��������؎Ɂ���CCt��
 �F��Cc~C�h CC7C�@�O��J���&C~ ���FE"�Bbh�Ga.F�/A��@�� ������F��C&� �� p  	� p yT �w 4 #����u�p60��{ ���&�@b�g�y���� D�Bh OBb|J�H��N�jkN�OODOyIH.���D�J��/�p�{	 
#jii�8$�F�
(?N�
O6kL�݃*+�tBh ~O&�I(OCv��fI��p.O�<�k�{� j)i8�!�jk��ii88B�JF8b!
�jN��
'O
'G`.F�/�H���~�> < U�z�w ��&z��| H��#bh�#��/��!#�##Ch�#|0�#d#�6##C�b(��h&��"ѥj��bh���&��| ��b!(�hF.4�� .@���&J.

���&��)⸕ [	��"�b!�� ��kߗ� �����;v  �  �  �  ��� v�    P     P P��e��z0�   0, 3, 18 0, 18 1  VE NT UR ED OM  G IV ES  T RI BU TE  T O  YO U,  [ A] DV EN TU RE R  [G ]R AN DM AS TE R!    ��{%�%
.

�r�%r �Ћ ��"�b�t)܀����=���ky� �� ps �+��@�6#G <@ d�2�%     �H� (�#�   � �   � �   � �   � �   � �   � ����8K��[���  �J�8� ��#���
�            �    �                                                                                           3�~$@.�(/�8���%�*@H��8�J8�k&.�%����'#"&?��+D.+&b&�%.%�k� �*%b@H��%&b&�$ N*�J+��&a.&n%a.%�k�@�,+"+n/&"&n.%"%�k� ������&� ��P�#[boڂ��o#?#�#O���J? ��           �L,�υ�	����[�)�9��	�Y��i��i:�y��y��yE�i��t�y���� R�SRQ��� 0�D�8�8E ��T��C NT(��C N ER���CR`ob�R1��D�8FN`� 0� R��OA�R��D	�` l.�σG� � 8�R1�� � �i � *j�W���|���+ �FF&D.�f�� �����
&

C  /�
���w=@&A�nqi0tiu0� ��^t)kT�%�'&�'0[b�ui(^�t0�ҵJ^t)e�&�F.���.w�	��Jq�����kk^�     Rڈ \�  �  d* �o�A� ����  � v� X v �      �����A�~
 Ӈ  ��B�¨�Ӄ������Ą�D��D��D ���b ���n��&�����b��f�9 ��&�� ��b����&��0��&��3��@!�惃4��@��o��F���/��"J������݇�D �慢�/���� .��X���ƪ����V�������ݠ��������O��L���8�}                                                                                                                                                                                                ?޷��� �&��6��� �d��'?�� �b��{ɩ|Z$&#�&&bȠ�%+f�/�?�#�&�&�#�#n��cJ� O�����O� ���{�"��n�㶯j&#&%)�k&/z�#?{z�#�:�/���i8�����&�J�����n�ss"��&k�? �v�� �v �� � �L̈\�c��z�F.@�w��&/�D�}"�@"�,��@��w##T.#""#n��/h#�6#O�#��w����&�&z��| (�����&�@.?��D����)ɩl��*w�֌��љl��+ �J�!�,��b�@P��\�މ���k��bX�Uޕ��q��`������_ݛ҉<���(��ۋ&z#�)�l�+� ��ϡ�w@!#&��6J.r���&��!���'#!&?��J ��|J��c�%b ��&�/��?�# &���,��{|����?�������������Հ�$�"�?��۫���  ���w��{HIݟ ��޷�	�֖�?���һ�ɤ���U�\͜@�Y���⃋l�/##�?$�-b�$��w�Z�(#�!�$ .H��a��?�-$&?�Y��J�Y�#�b�$f���##c#O�-�#.6#O�#�/�l�����'(f)�n�j���"�rH �F���'?�����+�]?�##c$#d���##c%#d��#&6?#�$#'#�J�#�%#'#O�&�#?{�c���@L�                     p��$�$bi������$�$�f,%b�$��.�/�h,&&�%&%.���+�/&�J%%BH���+��Oc%��$��/$(/? �a?�Z�>�.b����۔/D./.b.�+%b���c۔ -�������-/b ��+�k/./o�,�&,&%��.�,b,�+.+-d�ܫ��H�/)�I�$&��������!$�$.ba.�&�+/b�����&�E�%."����,&�%�%�%."%��&�&�,�J�/�,/�@�&.,/b��a�&n,q.%/�%��+�@��@&��%�&.&$d %��%��&��!�%@n.%"��% n++&�%�(&�%�h&a.&o ��               ٵ����/)݋/�a/�.�a.������.��?�%�/�$�a-�`��!��@����(a-�$]i�?��@/���a�����?�� *�.@.H�.�/./-d *��,�k�%�(&�(+����%� ��&�/���YȚ$+f���%&f� �                                               +,f���/�                                                                                                                                                                                              v
                                                                                                                                                                                                