����     E    ?4:2
$ 6(  .,
4<'> 8   -
<='>! 8   -.,  w=8>6(x A 0< 2    2". $
%' +".*  $11?  $ ?$)#?
8 <> ) +0>5 ? ?                                                                                                                                                                                                 	� �@ٔ�MA�':�!�    �                      �                        �    h��     ~   ����� S0@ ��  ���$���K	g⪫f� v1[��V�U�� �HWM?t�)��T�� �J ������ޠ ����� ?  
 D B��D���)~}��n|��{iz)5�� �B�{��1�{A����L�; � �yx� �F���� ����w���� �v0 u��K �&� �tʘ�Ȫ�����K �@������+ �@������+��F.������r��/��朂� bx�/�|��خ wb�n��u���P���?���������X0��� 0 �/s~��u�s ��
>

�����r���K w (��qw q&u,�(/������)�p���o�n �p���r��"淑���;M� �E@u����B3R�8G  y����� 5`���PŃ��I	�� @y���o��R1��D�8S�ny�aih �    � �� �}�m����C`��LS! m	�� �C@`�XC��1 m	O�� �
� E���`TpBR�� m	�PBV�����mI�PBV�����@��Dm˔P(V�O m��ɄSV��m�NSDV�m���OB�m9# u�m���� 5��SRV�C@!y����r�uk���2�ހ��� l	������k�� otI��/�k�O�����x ��c�(O�������J�6�� �.���m���� `[��	��DDO�@6y �.���m���� `[��	��ETm!�3 y �,�t��@����,fj �i�F.��j�k��+ҀHMw?�A)�E��@��JH`� "}& �hz��qO�}O1v�sO�O�O�eO�kO��O� @b��/����t�p�����r���j(/�h�gb���ֈz��rO�}O1 gb����j(/�h��jg�(r����( Gr�� ��vu� ��oi�"b����&,!�ʀ�� h	&rf�	�(e����ɥ��%� � �|d�c�z��E `   b|�da���z� �( `b|�da�z)�E��G���       �b��`��_)y|�da�z)�B��������    b|d�aј�/x�z�#�T `b ���ti(����/x��|�(����/�^��n|�t(����(����/x���k����� ���_:;�F@� �,�t]����,fj �i�F.D./i����k,� ��+ \	�\i��b��&��/���DXf��
     [�� ����&��&��l�    [�&�&���&�"�l6
.w��n�%6%"&&c�&�&.�� �'&� ���&��J��J� ����~�%�H+� ��P���2�y�m���� `[T�8�OA y[m`��� `[T� 0ym�`��� 5`T�ƃ y�r���� ��i  �����/�m���� 5`o��R1��Dy��y���y�(/!�#�b�#��y�����/�� #���(#�Jy�(�!#���(#�Jy����w�p��fـfɔbFx�[$Z��K��y���
�
j��y� ��/
.
j���-�����b
�Z !w�F���&��"��y � +�x�Y(�x/�/X �i�W��.�hV!��hV!�b!�(�����&�.&ܬ��/�/�F�.c�.�z ..�"���.j0{�/�.�
�w�H(�����$�H�� ������� l�y�b(��Ț�(/�!���b�y���(y�(��!������y���   @���y���b���(/�!���b�y� .�i ��@������*b�������(y���y� � � ����b���� �U�T+ ���ڨ/SR�� �@��T���i ��@��T�y�lv6� (A �Dmi��� 5`o��R1��D�!&��&.o���!�Jy ��������ͪ������m�W�N	!�@:�m�ԣ@��m�LC RQ��D �
m�RT`Ra��D �
m��@:�m�C�� 1�3	X��3��@@��m�MN"�R��D �
m��@:�@��"�������yº� �� � �����m��EÃ��#) P�m�A� �PR0`R��D �m	�G1LN�PO�# �m`��R1TO��3 EV MRMAN ym���� `[T� 0y �� ���H������ ���b���ĲT �� �@��TջK)����&�J��' ��&~a.i�6��ik9i�2� �C ��Cȏ( �'|)�dt�zF��`��S�� �x��|t�(x���/�k���f�	&	`?�����	�"�	��	c��f	$6+b*\i��/�*�$c(��$QI�$�$�i$��yl�P)�)(/PO�)|i����m��N�Rנ3TBT%`��A��P  �   y �+�N|�*�k�����*$*B�j ��$&� �U; ���B �q�S� '(����i�� N&� �&)�/��((c@�☝�((?�)����(�*m���� `[��	��D�A� 0y��m���� `[��45N�R y ���i��� N�m���� `[N�Rנ3��TO�#�8	�$�#�4y)����"P�U���k꠹��D��E�S����7RK�"��/� @�i���K�� �K�����I�� �Y�T�@�	                        
B �       ���	 �       I
 P�*2�1 �       +������ �%7�X��]�b'�v �p��             )
�2��8��A�� �            �q��? �F�W��� �� �  ��  � ָ� ��� ��  � �� �ψ�ň � �� �  �� ��  � ��  � �� �Ԉ�ψ� ��� �� � ��� �� �Έ�و � �� �Ɉ�Έ � �� �Ԉ� ��� ���Ԉ� ��� ��  � �� �  �� ��  � �ň� ���� ��� �� �  �� �  ����	�D� �	�� �� ���?�)�z��1��� �      M��m���� FP����LX� y &Ȩ�m���� `[� 5�.N�R y +�x�l�b�����(� ���FD�+.��|� ���DD�+.��ˀm���� ��OB�3RQ y L�K����q�n�@ ��J� �	+F.����{ �	+F.�!�� �WJ�� �W+������'� ��)�z��1��1��1��- �   M����/I+������'� �Wt�(���/t�x��+������)H��@ I���b�&+�/���&� �'�'���&7�'�������? �� �2Q�� ���Ю h�����
 W	H��@�I��+bD��&7�m���� 5`U��HA�M�`��Ճ4@y W	J�� ���4(��!�l��D.����k�!.���� �{��|��� �               $11?  $ ?$)#?
8 <> ) +0>5 � �J�� �H���� I��+b����'� ��H��� �I�&@>u�/I+��G��'� ��J�� ��ۈF �E�n"�E�H����I�cv�b�!.s�{ +�x��^�(��,b�x�D �i�� ��)�z��1��1��m��m �      Mۻ t	��/�|��k��C�������� �m��L#� �Q y+ ���&��(�.�枎J� ��FC��       ���B	�c�!N!�c!�	C�/�!�����	B� �+�/xY��,b�x�t�(/����x�&�/��"@��i���"�b���Y�,�/�t��x��'������~��~i}&�~'�孠��������O��L���C��� +�x���*�bQ��*��bQx���"��{ )z��1��1��1��)��)��) �      M�� �+�/xJ�� ��+���{m��N�Rנ3��ă@y +�x��^��(/������ր����ր���� ���d��6��C(����&��7��D� �   ����������������������n���� lg��� �� �� �� �� �� �  �hBL�D���a����/>���bń��'��'}'�P � ���&����� Ь����i@  N��&��'�@�  �N�� �
��������������������������������������������������������������������������������