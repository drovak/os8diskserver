���� @ �@ � @ ��	<(/2	',   *"5< 498
+/     o4 ?0:, ?= ?&?< #-'9?p 6:   ;1*>3;/.:=6-61  -;1   81+1  <12302  
<1203;  
<11,62*;  <?34   -;>4  
	-;><  	-                                                                                                                                                                                                 ��/����1��!��]�1�B_(/ I                    E                         3   8     @=          ` e       I� �m�TA�Qn*e�RS�"���B"�  �
 @/ـ���B(��X')��� X"'ӛ�t� \'e�'� Y�Zb^b�t����������?�ڣ��ǉ����D��� ���H?�����'��<�|�(?��'�(?��'���� �
�����r��r�|���� �
���� �
����r���ˁ����s�����D��Dʁ��z��ˁ1�-����E�D����D���4��*!�� �>_?0P3������N%ņN�PO  	��L��	5� 0��P3Ne�O B4CSO�#N�PO  ���N5�O ��	�S Ւ@�	5� 0 ����2T  P � ��(��b�b

bb�ن&[�& 
� `�6�' ��tׁ�� �/�i	a>�/�	�a���	a>�/��� � �~ �� �                                                                                                                                                                                                ��,��|�>��l��;   �|�������������� ������ ��.���� �    P     @ `     � @     �^    6 p�M� � k ��BA�խ�PlO�6�ѝ#MLt�eS�Su_������|uS~�@�� č �� �                       ��� ���D�Ϣ���У��A.�����ۈ�� П����&��&��&�Ϥ����������� �������c�J
��

��J��0��d��0(���(/���(���(/��(������ ��������&���(�����  �Σ� �Z.
����C��d��d� ��           �� ����� c�g�� Ѐ�N������ m� ��1N� �A1�2� �1��� ��1/l�ͻ �?� ��{K� ��{+� �Q{+7|� n
{�r �`�>��� e� �&�>�m̱ Ѐ�.� ��q�s�� �.�� S�����} ���>w{�w�� ���; �:�,7?� p���r�� �5�0�� ��7�2 ����� �B,+0 ��w^| �                                                                                   ~���	�#1$                                                            �! �                  	   @ٔ�@    I � �   � �                                  �    ���D P                      E           �  w������ ��@`�ȧ`Y��+�u ��TOc?p֙t�3 �Q�"id�8��4  h4߇�8X�,���əL�(��M'IO��a�☀�~�&�ə����b�bI�b"�l��L�/�N�"t�N� �j&� �"t����/� ��/���j!.�"&}&|6�X{��*�6�bz*�zy�B��!~iKx9�w���v��~��"4�u�!xi�w�`��vC��z)tu�!yi�&� ��#�%�=��x��� ��d�c�R�R$��sɒ$����u��L�?�� ?�~� ri!6⠲��z)rz�&5�/~D�5�j5F�z)�+f�"&}&7"�J�5�{ɚ�z)*z)tw�������
&${i�*�q$�p���w����$q)vt��z)r!�$$b!z�
&
z9$�Jto�x���z)t~��t10 X/���&  n	X��vm�p������z9qw�������yߖ7�w���(/��(����/�ߢ���lF����nW���$"b%ui%q)$q)F�*ߔJ ��@���~�tKox��w���� ���z)������r(��F�u��z��zF�zw�������� �r������z)t{��z�*z)��#zn�W���x��� &�2T��O on�Y��v��nW�����t�v��RniX��v��nT��v��n�T��n+��n�T����zl�z��zn�W��wt���/�~�t r	ri"�kn.�mk�A@  t�n;�mw��o�v��z)tz�jz)��� n	;m������¨����fffi�h$�����$�*&&&�.��}������gn�2m�k �  tg�kB�@ tn�(m�gk�C@  ��Jtkgw�m�����КnQ��l����� ������'�k� 0�t
��l�G�(?�ۦ���#r#r!#�
É�#�J�w�t��nQ���o��۱j~ϐt �k �� �t��z"�!H�zf�te�F�$�f �e$�n�;m�vm��z)t-�. I���� H!�/��������&��&H�,��|��K   �(/����i��� �
��D�d��� n<�mw����m���z)����������-  ������1  �
�&''?'�'>'�'�'A'B'C'J'K'���  �z)5tK w	�c�(����/����Kn4�mk�E@ �t���! $�� �gn�;m�nX���=fb���%Á�����%;&�7b<pi�ê=(/�!�=bc$c%�l%�2%%t%7%'�;�<r$r�|=�Jwt���/�~�StK~L�t=�b���%����;�?���<q);q)�%����7�ށ,q%�q�� �%;&�;�
�n
;6
72<
cށl����� �� �� �� ~t �� �� T�� 07i�l�%�%Á�����
&$%b9�w����/�o��7����,q)$pI����8�
&$!.$�lZ%ᨁ�9969$2�������9��
�:8b�7�7�l9>		c	c	c�la:�8�(8�n99&$�J��K�$⠁��
�7�j �&����@��:.:d�:��9� 9��?��@��X�vm�{���z)f$�5�JnT�t{��*�z$��t��+��z)� �+�/�~�It+y��l�$�$����$���$�|u��x8�H@.��/t`�zz�t~��tKg{�m�ml�FniCm�5�H�F�q*�q�tk z	Fz)vԛ�z)nT��v��w��ݢ���vԛ��Bzԛoz��z)�~�t~��t3�)� _ ���('  
#f�D6��CE�d֚lG�GG$q#��G�E��D� G�DG'�w���� ���@�8�&%�k&���G��Z�GG7G%BGs G�G'8'@'%r!%�Éǁ%��w�������o���~���~��~���J~������������n�;m�vm��z)tn�2m�gk�D@  ��Jtk �*�T �0X !����"����(?����bl�a>�à�����e������Á������:�7�'w��&��Éǁ���e@�����a�☝��~���K    ���d��4��b�!b������(����	&��&�	�a���?�¤؝�����6���r��r	g�	É���J���z5�t+�-���  �qq�w��(/���(����/��������qz��z)����/���q���q)�o���l_�^�����].��\�]/��\�w����/�o�]0��\�w�� /�y�^���nT���$b%b ^i���n�W��&&&$&%& &d�]i1�\~��[~O�[����fX��8��'�B
	$���U� f	�Z� ��f��Z�/�o��Y�e�a(��`�$�b)�b��b%%g)F��%)y%%7%�D�~�[+�&l\� $��f��e� u	v��w����/�~�Mr9���r$�$o�r(���$$czȚr�$$k w	���H���@/�����Koԛ��/���� ���6�wI����� �PH���n`�?�'W����~Ӕ[$�z$�zw�X�� ��R�"���$�L�$!���$�2$�|r�q�v[�p�����zr�zw�X���$�z$�z��^͚����a�:8bW8�%B�/���]0��q�p����@8"@�j �G�<�����l���������8%d ��� ���4�������� ������*3S��U �}�X� /������ ����*� /�w���������*o����� ����*������n�R���Á�� 	����l�<(���/����<�?������J~Г[�r(���!>�?��q�q�CzĚ "ܠ�"�k�C� �"q)q)� ��"(��������+���lǶ���V��� �� "���"�k�2(����$� ��! ���z)��4z����4��{ ��n&��; 	�n�R���"(����/�����K ��zl�$$bzw�������$�LZ$��!"���$�0�V�/�$��$'���z��r�q�v�p����zr�z�o���~�O�;~Ӕr���~���J   X?� �` �a.�/�!�~�t �w��eF�wi���e�� �f�h���(���F.��h���h�F���h���h�F��]i2��*F�*����@>/ρ|���~L�� �wϛ�@/���H����$�o��{��s�����x����z*�zt�~S�t �&!�� �~ �U; �,��
�F0�� �@ @ � � @         	  
        �""&���k @"n"n"n"n"n"�k��4(��WĚu')�)���I�  � �
��'�b(lb�v�-�)b���"P�U���k꠹��D��E�S����7RK�"�&�p2 �	!.&��&.��Ȑ���)�����.��b��.��b�湷����b�b�b�b�bf���         ����X*�3��#(?���%!>��/�%���J�v)T�&#!>��?������ᠮ# 0����#�##s�%&�%'�!.%�"�S���b��f��&C &~�*�qO�? �F�W� '&ffff�wi�ָ (i��U�(Bbbbbb�i�����ff�&���&�/�w���� ��y���u�o(�����&�u��o(�����Ί߀��,F�њ�&�����/��� �(�� ��o�� �wߛ�H.���'�J��o�� �vt��z)t"��<�SX3�G�
�R*� ,i��U,D.D,�D⁑�w��� �������,!.,�hV'�^^7� ��&�&��(�!,�@��!,���*,�b��b,b(��H,�����cccccf��ɳ���* H�.b�.b�.dG� D�.b�.b�.�k* ��3R�VJ� &�&�&�&�&�&��&fff���H��.��b��.��b�����J&���         (/(/(/(/(/�/�ڮ /��(�(�(�(���������j�k ���b�@n��q������d�ث    $���fI����K��� �����
3*��į �	����&f�����i��F���u����t�����i����7��J g	�z)�b����z �%z)7z)�%������wҚ�(/���������cz$����zw����(����/�w�t�����~�t~�t f	�Z� ��f؛Z�/�o��Y���K jz��z�z�z�z�6  �T� 5*	���w��� /�^������nT��^����n�W���� ����*�(/�������Z�b��f�o�^������$&jz)$!.z��w��� /�a�(�� $��)&f%��&)֚eF�)i�e�'%�J�V%�������'�'�'���o���z)az��4�  �j�8����$!�`�/��X��                                                                                                                                                                                                �$&Q&�ɀ������'$�J� �$t�P���/�O���/�����ǁ�̸	���ì�t��D�������ɀ������`�=�����w����������������������������������������̉�����������ō�������������������������������ŉ��������ҍ������ɚ��(���'IO��a�☀�~���������&&&�I&�"&�ɘ������'"�J� &� �"t����/�������� �"���&��!��"}byi�&�Á �٤�&�Á$�$$�s�!$����Á����u��L�< ��u��dӐ�����`�=�����x��w����&�����ni2���C��ǁ��l�AAb$�
&%�l�"$�|nX����l�$�$à���$'� �$q)%pIͥ�%�,%r!%�B&�
�
c�ǁ%��t�C�/t~�tKn?��d�C�b�l�<(t�$�b$�zT �                                    J   AB                                                                                                                                                                                                 