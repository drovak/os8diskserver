����   	 	:   	      	           @  %            .                                                                     '$)  +  2A ? ?0,=                                                                                                                                                                                                �+&@ٔ�MA�� ���L �   �� �� ������ e         �                                           ��       '��� ��3 �D2�_���? ���� �� ��� ��U$�@� wQ�7�C�E� Q� P����w �O�����ڈ��y�0 ��yx2z}��$�w��v)̑�&!̕?�?!.� /����@&���@�n$wiuv)����&!̭?�?�"(���?�tH/���H��s��w�?t"b�F&FF6FF��w�|���~��v �����b�b	�b/c	/t����z){ �}����|u |)���� ��G��~ ـ�� s��~|����z)�})��{�� ��� � �  �� � (��vQ�x"z}����vK����v�uv)Pr�55bq��5x"z}�uv)Vr�66b!5�(���6�q7�89f:pion��v�8��vܛ���pJus �խHt�c�%\�� �AP�CrR� 0                   @�� ��&!̅?�?m t(/�s�?� (���v�뀲m�&�w��?�l���v�� ��v� ���v-��� ��@f�)&v��uv)�r�6vil Ԁ6�xz)}��)7&7�?�6��z)}�́�~ � �� 7ck7D>(.9���6z)9})����7@?澪 ���� ��?`?`��؇�� �"R(/ �?�?� �(/܀�?&,!��w?�!A�(���?��!�(/���?!.�(/���?� !��(�����(.�( d���))&�)"H���� �K�)�H��) d�����~P�~�ʚ~s�͚ �K�@ʈUi }  e� ��*�� �  D. b ��l�Ub!�l!t=��!�p�� Eb�<1� U�� )�"H���H/�����)��������������)���6.*�i��7�0���!�"!"b�"&�&��)!�	( ����)Ԁ�����؛�7��6)q��5&����9�/�8�I�� & 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3� �0���� w��p����v�@u�vV�r6�6q)�v)]���&!̑���P�%�w���j)v���� j�v�����jv����� .jv�Ā��j)v㜀�� j�v���j�v��j�v'��v)�&�*iih�v9�&%B ��g �.<f$.@�$�n/�l.<'</Dہ�9:fon��9�:fi�n��ѫA�� �
��)��&�@��QD��
ӲL'���v�Lu�v^�r6��6�qڞ!/�.;f9:f�;ǁ;�/�J�e��2�6:"�3&94&d9�:�n��v8����vU�uv)er�66bxz)}6�q9�:ei�2�c6":3&94&ds�9O:nI�g�����ݢ�!|�ԫ�����d��6� �   �ۢ�݂��d͊���  ��� ���J� ��w)  J
�
��(��H����v�_u�vC�r5�5q)uv)Jr�66bq��5x"z}�6x"z}�78f9:fpf��È�g� m0ei�9�l

�x2&9b �a�`6":3&94&ds�9�J: N0�J� ��3�����4!.�(/��N� ����/xb<;f�;�!<� ���;�</D؁��� 	                     � _����/viku�vg�r6�6x"z}�vu����|�"A��4�6�z)4})��{k� ���|�!./A@��4�6�z)4})��{k� ��4(/���s�/�J���/vi~��|�6"z}�Ԛ{k� ��|���4�6�z)4})�{k� ���"(���Js/�����/&�� 6_-�_v���&�6�z)|��}��{�k �|�!.�a��4n6"z4�}��{�k ���s�/�Jg��v�����v�xv�#u�vV�r6�9:f�:�9�_

�|�`:"6z)9})Κ{-�-k  ���|�^:"6z)9})ޚ{-�-k  ��9�J::B(���]�9 /�g�\v�+g�        � P6� �m0&�7�l

�27bb�a`"58"37b4di7�J�8�80d��� �m0&e��9l 

�2�9b �a��6":3&94&ds�9�J:�J0�J� ���,�n~��2|)3z)4})ʚ{-�-� (���Ú� ��:���9_ 
�
���  		    	     �x ���!�>>b�(/ǀ�>�"(���>��(/��(���>��(/���>� �>&>�"(���>��(/���>�"(������$��$�v�����΀о[���[�����   5454   5 .   1'  0'  525�X���� �@ ����� ��  ��$��о[u�v[�h�*&ih�Zvd�3.�4�_

�*iiYv)~4��*;� @�
*�*iiYv)~;��*iw�h�Zv)n5�l�*iiYv)~��;*6�i�h�Zv)v6�l�*iiYv)~��<�<*iiw[�s���� 	     	  �  0 �m&m+&*.*�n*.*�*� (��>f>X"W+����(/��������V�* @  %            .                                                                     '$)  +  2A ? ?0,=    ��=6��B��n=>U>���=U0>�h=�J �>(/�_��>��/�>&>!.X(/����j@/���V$���>�(>!.�(/��� �A�(�(� �>$b@���H���>�&!�ˀ����>�-��ڀ�� �$.P�$�k ��!>�nVW)��J��K �                            @�  �$.���[�uv)Jh����!�"!"b�"&�&�v)!h	ZvS�-*&ih�ZvV�3*&ih�ZvY�4*&iw�[,�@���-��(Հ�3� �z)�~�P�~}�Ț�~�̚,�K3� �3&������ w	v�v�v �v-�v@�vL�vU�v_�vk�vx�ww����:,S���� �-�?`��0�� �[w�v��v��v��vݙv��v�v&�v=�vV�vm�v��v��v��vؚv���[��[� ���bŽb�F����!�b�F���""�k   �"     @���"����������`�0��p�8�������� ��ڴ� ���� �� ���� �� ����                           ����NTR�.�S��� H��AM  n�R�	��E�8��AM  ��A LG�N1 Tǁ4@�<T�`��D�TD��EC�8��AM  .�S�"φDN!�S n�S�"��T��MS���$D�  �Ѓ`�`PR0S�#S� .^ÀLRTN��KS n�S�"�����4 0�C���AM0y � *L) ҳ(��C�iC���	�S�V@I�`��S@Q�TRSQ� �  � �N %#���5TXVC`   �  � �  � �N %	�4���C�SC��`Q�TNL     � �  �  ���C���M��I� �Q�E@   �  �  �  ��R1T���T�����@R   �  �΃�SB �  �  ���ԁD �D�0O�#  �  �΃�SC �  �  �B� U΃T�#    � �8�`1�8� H ���T�EL�C	� 0  �  ����@�OK  �  ��T2���N2��    �  �  �  �  �  � ���R@ TN	%� 0LG�N1 �QTRS� �TO�# �1�Dǁ4S18s��@6  �  ���C�-�4  �  �  ���@	�0T`V@   � Ҁ(���HT`  �  � ׄT� A�RNR�LG�#N   �  ��ң;��R1S�`�  �D��`1XX �UDN�    � `�  �  �  �  �  � ���Q�E�SS �TRN�! �T(�8�$�R��ϔNE% A�I� SPL���HKS1 �I�3�T��RN����AS���@PR0`NT�.�U��: PN$ NUT�.�5TX�:5 �8�1XS? ��0���X��0S�:Q �KS S@`@�KAS� TS`���KS S@`��D L�G�#NTR�O�N U�C�N(��E����38 IÕ5��E�UK �DDP8
SNQ @[ŖD�M0 D@��$E�3@	��HA LG�N1 @[�5� @PT� @ ����3Ѓ`�cXM`	�  D��� `[��D�0 �K�LBTO�5�HS�%���EI��4 ��		SXC��  ՃTU����4XN`!NB�T R��D��0�DAR�N�!���	�����4 8`�ǁ4`B0� 5�T@��	���C���T@�= @�X�	H�4ǀ>�,��@� CD= �����,Q@_� NTRT�}   �RQ�`<�P5����4S�`6���ER����P3�[̓MAN �� E�� u�u �ER����P3�[V�R� �� E�� ��� �ER� ��P3�[̓MAN �8VR� AϓT �P� Htt� RQ�`=�P5��R1�51Ӊ��0Ӊ r�r �ER����P3�[�R�0X���18� ���� RQ��=�P5��18� ���� RQ� >�P5��08� �00� 	�H�`1- �L ER�����$D`V@�O�5`��@��`1V@!��T�:5 ���A��: P�C�DՃ	�S  � N�T ( �L h �A 8C � P	��	  @B�DRD0 �  5�@P 0��D��@ R�C ��  �  P�  �����������������ҕR0@�a�A� @A�4 P � CA@6��# � 0U�� @�DM���C�P��C�BSR �BR1  y ����� ��
���TՀCO�3