����  � @�%2$2#2"/!q!8 '%$*#"*4(!4+"$ ?0?> ?7 8?20   8r   3<": ?*
<>.   0: 2?8 
22:/>  : ? *-
230
.0
/11*#0*!2?*22:'=.?9                                                                                                                                                                                                     
    �    ���L �                               ��3Z�"�n_�# "DS �gf-f����J�j�� � B   B �@       �#D>�D��D U:�U��U�.�8�� E ������J �̌v��? ���   8      n�f�� �AAo � � Af �(��Q�(��DQ�A��A�C(���X�  �A�A � � �A��� .n n �� ��  � �  ��  � �  ��������������<��JO=��� �oD����oC����oE��������  �਷� ��h ��h �  n�ӈ �  n�ӈ �  n�ӈ&⛄ �&�&��� ������ � �� �?'	 >�'ě @�� ��B�	 n	(����� ?�'ך @�� �>'	ӄ�oM����oL���oN�������&ћ� �     ���*
)��� � � �.i�/����B�
)i��� � �o �.��/�����+
)��� � � �.i�/����,�
)i��� �
 �o �.Ě/�����-
���� � � �.i�/���� 33 0   @ �   $  � ��" �  � �  ��� � 呂�� ��ࠤ� ��K��K�koD����oC����oE������)���� ��� � � 0i1 � � 0i1 � � 0i1&�⸻ &	 &	����k  A@    ��        �  � @   @ �H/ �f 
� n
(� � � � � � �o��  �A�� ����)v n
(�� 
�  n  �� � � A � � ������k�
�  nN  �� 
� �N��koM����oL���oN����� ��&�غs)p&(?���A�o �4i)3�&���2�r�� 71� ��(f�k ��(f�k ��(f�k ��(f�k ��(f�k 1�BS�d��6����b����/��㨠��D������>�*�!&�!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0�H> ��	6�	Cb

�
���(� ��(���H��>�* ��� ����*�')�?������  &!�ʀ��@ �       B	�>�bWr�c�t�ʫM������ݢ�!|�ԫ�����d��6� �   �ۢ�݂��d͊���  ��� ���d�� �v �J
�
��(��H����R�lf���9^r:�r _b`b�n�b�n: � 4� �5�67����Sl&l���9�^:'_ &a&�&�:�  �4� 5�6�7���T�llk�_�9�r:jr �b�n9 � 4� �5�67�ǀ�Ul&l�0ID#��&" . ���a!"  ���&  . ���������3����9^r:br ab�b�n: � 4� �5�67��V�llk���c:'_ &_&i&�&�9� :�  �4� 5�6�7���W�llk���d:'_&i&�&� �:�  �4� 5�6�7�X�llk��D�B$ . ���a#"  ���&" . ���a!"  ���&  . ����e:'_&i&�&��  � :�  �4� 5�6�7���Y�llk���_ &_&`&�&�f�:�~: � � 5�6�7���Z�llk���9_r ab�b�ng:'�:�  �4� 5�6�7Ú�[�llk-UH ^ ���a#"  ���&" . ���a!"  ���&  . ����h:'_&i&�&�� :�  �4� 5�6�7���\�llk���_ &a&�&�k�:�~: � 4� �5�67����]l&l���_�:jr �b�n: � 4� �5�67��̫��e��U!��� !����&���� ^ � !.ݠ/ �!π��b���� ^ � !.�/�� o��� �  �� �  ����� �o � �� �oC����l/� ��������'�o�D(���� �oE�������� �&��)��` 0i1���o b!��� !����&��Q�U o �!��� !����&�d�g o�!�� � !.5�/��� n ���T.T .�����o�M��o�L�o�N���� &yڇ�Rl&l �bz�.�ഷ"�b

�
z�b
��&&��� �  �0�������!����"���& �  � ��o� !����&����f � !.�/ �!π��l������ o �!����;��!�##"!!"!#"#!"!#"!#"#!"!#"##"!#"!!"!#"# .4� ��7�����' poD����&u�&Κ�!�1i�#�1i�� n 01�&�oC��������� �!.��!!b!#�@�����& �$$b %��� ��1. � ���1 � ���?�.���?�. ����!�� n! � nC� �� �� ��� � ��� ���j���� �������/4�3��7��������/4�3��7�����o�7����� �� � n��  �� ��� �� � n��  ����k  � n�  �� ��� ��K             &�!��� �	���1 . ���� o	D��&��&����1 ��1 ��1 �1&��o�C�����/� �LG�2                                  ��"� P�D ���2 @����ͻ                                                                   ���w�$� ��!.������������ � 4�#�/�$�b 2i�7����$ /�!��������������  �4#� ��$& &2ܙ7��� � �                                                   �$� ��!.������������ � 4�# /�$�b 2i�7����$ /�!�

�

�

�

�

�

�

�

�

�

�

�

�

�  �4#� ��$& &2��7���JoM����oL���oN�������o{�H
�}oiG�����&	��� �!���д왴������&��و���}!.|�/����̲M�& ��  �|��~&�y��K"� `�y�y�?�|��~$����yè����� �~�lK� ��n|.!�ʐ/��"̔l��&��& ~ ~~ 0!~������~�J� ��~&�')~�J� �~�b'��'~��� |z?'� �{
?�'�i������x ��  o	D��&������� �oD����&�������* o	D��&������� �oD����&�����&oC�����/� � &	��$  !�0i1 � 0 �1&�ⴻ.8/��8���.� ���.�/ ���� ���<x/��<x/��x���.�x���<�/ ���<�/ ��.�� x��` �  � R��   � �ML%TD  � ��kLR�  ����R��� �  ���Ɂ  8 �ML%TD  � ��A�7ށt�`0  � �N  �  ���D�7 ���C`   ��� H  � ��G   � �SL�W��sGN"L   �CL� �  �R�  �  ���� �  �X�D  � C�LP� p� x �ML%TD�S� �QLD! �  �M�LTPDLS �LD � x �ML%TDR�S� �QLD! �  �M�LTPDXS �LD � x �ML%TD�S� �QLD! �  �M�LTPD�HS �LD � x �N`D0 �1HI� 1� x �N`D0 �2HI� 1� x �N`�4�E�HI �  �N�`� C�TI� 1� x �N`�4 5�HI �  �N�`��D�TI� 1��tA 1��tR�3 �� ށt��3 � �T�`R��D���N ���4�8M�`eN��  ������ �&� (����r��b�!��/����/������x�b����s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��s��{: ���D�E3: ���@	DA�0��0,�� � N�W�*ט����!w"� �� �� � 	p � ��8�ǰ� � �����Ȋ�/��� �����& �⁺�� ��������&�°�b��d��������&������� �       ��/�o���b������H
}�}|&���M�& �΃T�# ��T5���8A	�	8�R2C � ��A3�8N`!�R1�� �DM�P��HG1̴�8 �@P��o�F����x�����NQ҃��T �T`!҃��T �DT` ��R �D@T�`� ��� @��NQC��R  �T`!C��R  ���  \�C�D �H(�M�@P�-)��N���� �&!��"���� �=���(��Z�&;')��J�7�'v�&�,Q���K@�                                                                                                                                                                                                