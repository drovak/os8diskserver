����A � @�8'7/:: "8!62	5>(*5= 4+2/:  772	3: 22.7  1**q1     +  
 !?3>$! ' %���������                                                                                                                                                                                                                                              �� �      ��   ���G\��             v��        H   �� �   ��               	�6~� �o�������� }|F{ R���t��� � lHX��0�L ����?p �/��"!� ���s��?u`@ �3�L�������O�����            ���06{&�z&0y9�Jx�����t|�����F�����⺀�D ���Á(���,��|� ��(?����Á�ǉ�?c��� �'�c�(�J�'�� ��w�v���c��� ������F.������r��/��朂� by�/�|��خ xb�j�8���D��H�?���ut�����si�"�?��u����(/r��(����/�?�u��Jq(&p���(on)m"���l� ((b�k���f��fj&@.(/��i�&���-�bb@���-�Z!�!�-D�j��b--c��&�/�-#hz)-D�馬 �       cb(��z��/��t��A�e�s��(/&6s��&��s��G���s��"������/���b����"���gi#�
.f"�l6������p�%g�!�
����e�d���/��"�����k�"(���(/cB(+�j(/�����������b)� �{&�&�k   �"���� �o9"9�k�0�6���6QE� ��/���a�`���$��t�D���bF�F.�"�~d ��   ��6��c��d��6�!.�H.(���/&��@���<` 
 >����J��J٠/�/���تj///�/ /�/��F�.�d� �   |�||�||�||���    (���`_�a^"� �/F.D&]
&j&����� �	" .#�/�"�"F.bj& ..&�� ~& �d����j�
c�ǁġ��~�������!.��h��/\�m�/\�� b� � .f&�����(�/�[�7 D�`b f�����J��ˁ~�* `f0&/�n"!.kb00&/�I�l0(?�D�otZ'���߫�#`s�&�K��"`b88k9&6)�YX'1�b)&36) .Pn�-�)�"4)bW�&�4s9�&9J.V1!.3&�9�fb99&�/�9�`11�l9`0�@��/�`��/މ�9'11D���,r-��k���& ."(/�2�9�J�)�)@.'�/�2�D��U8&���"�6���9������   ��1��sbZ"n dg!�\¸\̸�b� /��/����b�o�?�(��������o[2�|�(��/\��&��&�!�\� �T �o`0!�bu��� .f&�.Á����K )W)"c!/����)�J�̋ )F��+ �^z)��J� ��!>@.��4��4������5����(f����p߀%�&���@@Du��"!.3fb0�jT?�u�o&(Cb�0d�0ÁH��y��Jjn)0J.V/����0�6o6�?Dc"6c`!�6�66c�n66&��&6��/��f^"16c���q(&�6����1z)�n��J3�J5�/r����JC�&T?�u�Cn)���f0"03d�ڪ���� �� �&�/��K�� U,� �!���&��&� ���p��S���/�w��O����F.�൵7�J.
�����r��d��J��(�����&��B��{    �
 � ���bŉlw�<�*�=���wÁ��*�H P�����&�����w�0���wv0w�z ������sP����� �� �=����&�~�~i�f�5��H ����  /���y)�z)�̈¨/�z)zz���!�����2(����)�*���ǁ�É�?'�'w�<±J�R�   �R�H P�ä������R�j `�x�   ~�~$�       p	����?(/j&���{��bz��j��h�J@ .?�k�� �� QzP�z� �	��@��D� H��� �� ���d��&��� ���J��/�����<����̈��������&��0J
��
.
�䪇�����C�(�R��(/����F� �� �    ���0 v�Z
d��6��F��� �@������z
�
��ہl� �� ��ݢ��&�w D��w ��b��b��k��O�~�$ `&!��������f� ��QP����7"2�� ���H#U� �M�� ���H#������ ����H�0�2�V�  0�&���J��	b9	�0b�����	&	�&	b9	b9�� O&�қ�\�� ��		c��b��/�ӫ�/�����PE)&� ��F5 �	�2b(���'��;��f`��/� �` �F�v��� ���j��F��"@����)��b�z��z)0�K    �i�Ģ���ġJc�'"(��o�/����/��E�N�/�Q�E��S���/�x�   �������i���Z�"�@n�.�X�R�"�cr��/�����s�fr��r��{   f �kFr� �e����U�ք�7|�^�i��jR*���>>�@��4V���)r��Vz�(����)�)!.�/���(�!��[�(���B
�b�b#~b
w#�J�k�i)(��h�&a.��6��bk�j����&_c9_�sQi�D ���_�r��& �ur� .&�jH)����&�J��' ��&~a.h�6��hj9h�2�� 0S�O�Cȏ(0k����*��<��?�w�������R
� 5 �
��,w�|����<�jb�l�<��t�D��������s����'�!'��Á��*���'���*�c�b�s�h�/��"c#c$cc	�h� ��<	�|�J�~� `F���
�� ��߁� �"�jCˣ�p�����OYr���He �� �	������<�������(���i��ʢ��rX�~��Á��(��R����G�����<���@����r��|�>��D�灊����X'��'_�'�T��|�������c��z� �큜'.����&��� ����'8� ���/�آ�'tс��`� �0��h�B����R�������ߣ����� �    8�   g� 0 �   ��   �*   ��   �*   ��  �*   ��  �*   2	�  :	�   \	H 0 {	~   �	�   �	L   �	H 0 �	D @ �	�   �	 0 �	~   �	�   �	�   �	T   �	 0 �	�   �	 0 3
*   3
�  [
�   �
�   �
�   �
�   �
�   �
 0 �
~   �
�   �
�  �
�   �
�   �
~   �
T   �
�   �   �   T   �   �   �  �   %H 0 )�   )�   +*   ,*   ,�  .*   0�   2*   2�  5�   8*   8�  I�   K�   N�  T 0 X~   [�   [�  ������3��      ,7"�!<& �`yο ��/��!�1 ҿ�� "�!�/�AӠ ��  ��Z�A��!z  ��  ��~ ��� �yI#���� � �+! ���#ҿ��"&��Z#L�!)�2� M4 �������}��#&��3��      �� #�!������&��� H1�O�!�S�+����M�!�� ,,"z  ������Pؿ�f�1�I�1[�"O�!yI#���+! ���#ҿ 2~�M4 ���1H�1D @ �FB�������� �E�i�E&�����k �	� ��{��B+Fh��'�¨����'��'��'�����r��r��|��� �"�F0�0���/��F ��b0
&�&
7�J."�l��0$��� �V'���"F.��',�b��{ ����� ���'�ҰF � @ /F�P$c2q��O�
?3C�wc��� �6���&���)����G���������Á�ϝ���b����!�	����"�!��b&����/��@��tǁ�� ���6��L��0Ơn��2��c��� �&t� �                                                       ފ��!"����� �#                                                                                                                                                                                                