����   ? ?(
 0 
,=,
&0 ?.6 !?:/ ( +=.(,0 &     ? ?<
 ?8  9�B B ���������                                                                                                                                                                                                                                                                        �P�@v&xş� @ ���G �                                                         ��`6�@P1��� τT�D��@��2W����00� $�_�� �l�� ��� !�_/� ��k�0n(��#Yp4 �# ]��@ ? �P���W� �9Q&��7�� �~޸/Q_��&�� f5�}�����A�!⨕�D|"Ȧ�ϭ�Q� !.�/� � �}ƚ �/��I�X����h*�/�h4�/(���jf�hA�/{&� ��z)yz)� �I��x���& �k ���d �}՘ �/�ޫ { H�Q���&�A?�� ��������썀 ���&��� ��y�( ���H/�|�@���{ @Q��A���j ��w������ �J �v�&�Ȩ ��(/���(u���+� ��6��F�>t(�ֶ�� �s�r�"�Մ�.���ԾJ��:      !��&��� �!#6%/#�0A!�#�?�!�##c�A#!t �J݅���� ���}�����s�&"b �� &�!&%6q'�%p ��-����o�������%p n�-������t���/��' Nt����%p ���" /���'!."�j�'"���D�"�mms!l�>�w���� mc!��!�b"�b@!� O��"�J� ��� ���:kYjw�� �������� � ? ��� �/���  '�_&�/�����r��z��'��'���ɼ" i	h�/�w�� �wg�R�/{�fe��� NR E���  �� �STU�ˀ�B3R����2�����剙AT� ES�q��)<�� 0�DT(E�dl��pz� ���A���8�0 �H��C�� �C���C��  P�) >� .d�()�b�*�4&5&/&�-����& .4b./b-/b0b%(f~+&,ci-/&.4&D�6�5�j56&6.&51&0-&%6�(�c.�6�k  0! f!@.m?� ���� .�� "��b �vib����C����%ab `b!qip0_�-^^�����t�]�/�ڮA�\0���"�JO�u:�1.&0-&(2b+�b,�b�ci!#& ~�	`n2
&  . &�)�!$� ��[��*�!$��"�`n	�b
�h� � �K-�/�#���K m"o	!>
�<���"�J$�J��]$"!����EkYiٖwْZ(/YX����� �xr}sw�w>w�w{0Wz)}�Z��b ��0t�JV��x9��IͿ7� U Tb!qi%�/GS�3(b � &@)�)��+��ǈ O��a ����p A�@*�*��,��ǈ� �!-�P@�-�k !-�!.A��� ��.b�!b..&� �vb�3 �   �v�b��-�/� �������g��l9E��w�R���J 	p�(�� @%.�Q�
� {�AW�z�H�$ �� � ���&������b��������&��C�d��6��L�D��������&�����Р�������'�H޿�������"(���d�!.��&P���"���퀟����Fޡ�(���/����� �� (�������F������J���PN��-�����      ��O �@�����D.8 �/��m����m����������&��/����P���̀���"���Š���c��?���J���ވ�ň�̸�̈����h����@�J�J.����ш̏��ވ� ���������� ����� � ���� !D���"��b �� �� .F�������f1D �  0      )����ɥ��%� }�V� Qr�� D&D*.D1BDFHDQ[Dg�D��D��D��DρD��A������"�� ����������8�:5 ���^L#� ��T� 5 � 5 L�1 �4��C� @��b�@n�u�N�*u��� �M�/|��� ���y����J���� ��|������J� ��fZ��_�صvw�����{�!���&(/�!���"��b�����<!�⨝�I�w ��!����H~�2�b��{	�!S �L VI�z �� � )���0���?�I�''�'}������~ /�ӂ�*���
� �    <aR��b��&�K"F�H���&�P.��/�󩀀�䈿���G���-��G+��   �����