���  $ �766%#%%  #% /  %    /767%#	%%  %#  +/2%% 	  #%  +T ')
)%				
%	*
76%   %%#%  				%%#%  *&*                                                                                                                                                                                                 c�v&xş��C ���G �                       8 ?  ���� �� �� ��  �# ���������� �����������@�� *+U��� 7VW ,
�C�� ��   &!�_"�]d���1](i;�0 8@ X` �� �H��=>U?zP
 d��  ���c��b

�
�菐(� � $ (��@/����>� ����*= /������&!̥������ ��  H�d��]���s!)��� ΀����!E⨴�!>:�/�<�]���� ��&H	&!>	�?�� ��K�?����� z (��~z ~)���R?�y	� 
��� X�� Q�A �:X��A3�8�1 �
X��A3�8�0��JX�� 	Q��T�`�3 X	� ��;�  .�b4�# �b 
��( �$"�b%�� n&
.

�$�.�5�� �       �� �    !�"���������&�!)����>�, l�i �ր�!��X��كC �U� ��Hߥ�����֊ �Fp"�-Zu�� �-�k��-.H����H�ǘ��Ӫ�⠒�XN�  H�X�A�4��� �X��D X�X��C� �X�	IS� 8�"�XiR��DS`0� Y	KҐ�� ��  M�"��k� �������
�� 4� N0 �Xc��X��T8 �Xc��X� Y�H.I�g�:b!I�(���,b!I�ȍ�/ .I�?�I�

�4�	I�J��⨊���3\ n\�~�\6�X�	��� Y	K͐�� �  �ʫ�K)�� �  �ҫ(KY�� �  �ګ KY�� ��  �
��KҐ�� �� ��  c�ȣ �F��!�zE�i�)����3y&�n&;!.�?�,�!��P�0 .�?P�"(�a�c/Q��J�J(/*""f@.>$ ����S�A"!�6&�3�@�OR������ .b7&W)X��1 �W�X��0��C�E���C݃c �YK��� �  Mk��-�m���XŔ?T �
$��� p3:�r"��&�bJ>r[Zy�JC&����� �J>r[rZi�ҲJ>r[Zy�J'@['ZݒJ>r[Zy�J�J'@['Z�J>r[Zy���C��h�J�bJ>r[Zy�Jɀ�J$8 N1R1 �V 0      ]� $� a� $�$ �$$�h 8 l 1 � �"����b�k�q.A�$ �l"����X�� E�TB���3�L@ Y	t"�D�d������J�J'q"��bT����n���� .[�rJ�}2��[����B['OJ'l�-�ސ��l�*  C ���c%��أ�e�ȴ��7�� \ � 0 ��\&� .��d��\�t�\�!����\�J   � 0             H��V�bZio�-�J'>['�[������![�J'T)���j �2�����[�����J'���B['NJ'�[�����ڀ5D   ?9�������Mȳ� 0��b

�
���% ��&�.(���&�% ��&�.(���&X �   � �0��dB� !��(�?0B��!@�������}R��_�����Ȁ�Ȩ&Lf'V) &[vrJZy!.v�?�j��[�wJ'[�?�L�!x���[�}H����j���O!��/�������2Ш���LҠ�� L���&&�ª(��! ��j>D�-vW9��WX����@؛� X�L% � ً�-wW9�L�WX�T�`Rc ���X�4	��ԃԃ� ��V�'�&�V)B&H	&GJ'Z�	t���X�` WX�� �B&H	&	W9X� ����M�� �� 0��7�J.
�O���r��d��J~�)�Ê��&��B��ry�/4@�~����� �=kR��b��b�@n�u�N�*u��� �M�/|��� ���y����J���� ��|������J� ��fZ��_�صvw�                                                                                                                                                                                                