����A �                                                                     A8 
 > 5?"?���������                                                                                                                                                                                                                                                                                     �,��v&xş    ���G �   �� �� ���                                 � �            ���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s�
��� �v��� ��/�?3�"2�������
 �	�������/����/����/����/����/����/���7� H7��H/�����y����/����/��j"F���e���#.B-�i���-����e����  `���O �� ?�!��� 
.

������ z (��!���/?A04�;8�V�� � �0�~)�&~��}�!|���{Á��/   � �"#f$%f&'f(zi�(/������z�������/����	&�&z�����	'�J��K� s -d8K @A� UC�0L ��Kn��Nm@����@�l�T� ��i��bi ��Xp@��u@ee�@ BP���s��!�Zf����� y	�b
�b	cb��/�
��J!.
�?������ �*O��yb	�l�<(��b

�
��	r�	�O����<���D�*���/��f f!�j � (���� ��+ z�����z������e�/z~��"���z��(���(/������~)���� � ? �"Zv��? A�!� ���K ��	F	(?�&�!�ʀ�� "��������!�h-D�.�-�he�K ��	F	(?�~�� �                                             �2@G�"o����""�j T F��{'�+��D. b ��p�Yb!�l!tF��!�zE�i�)�}��H/ ��/��������+�3&�6&�!>�76�F.�7"h��J
�
!&5 �  p�6����6466C�6��J
4�

�6�3�J�F.&���>&����B�/����)�) &�)�����4(���/�פ�ף  ku�D)t&(?���H�s �=m)<�&�� ��VU3 ���f �	��&��&�{�(��������[��*�&�&�����@V�Z��,{�|�,&��'��'�	&�	�(��/	c0	c1	c(��2�l��&��Á��   �
�|'�+&�&�*&����� @�β���� �
�5&���K�����@xiw�K8)���|ly���a��/�/�2��?� 6À0 R �6f�b3�c��r��r��{ ���x��hb����t�.�ଫ'��D�������;       +��,��  `�����b��d���w�K�ȓ�����;����װ�� �� �� �� ��  � �� �� �� �� ��  � �� Ġ �� ҍ �  ���   ������ ���"� $�U#  ��� �� �� �� �� č �  �� �� �� Р �� �� ��  � �� �� �  �� �� Ю �� �� �� �� �� �� �� �� �� �� �� Ӻ �� �� �� Р �� �� �� �� ҍ �� �� �� �� �� �� �� �� �  ��  �  � �� Ϡ �� �� �� �  �� �� �� �� �� ̍ �  < [ ?3 l [? 4l [ ?5 l [? 2l H J \   0� ��z���"�*�.�1/b0   ��%
��NB��A��C"΀����/ ��" �BU < ur��h��/�ⲺO��^"���d�*��~,�(/��kr����$t	c%� �)����ɥ��%� }�V�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                