���� d    	 	 	 	 */$0.1-&5&4:45&. /&8030-%  ^   ?98
<(*
8*"288
"2-8 
- 8-< 

.> *"
-*
28!;> . >=.  _=/
??A30                                                                                                                                                                                                 �+       �6�                            �
                        ��� �������� � �� ����y���ρ�����_���?�
� ��  3�![��*#�=�$�	g��f��b(���J�As�k�$s�&�� 1 &'V��` U9� �n�f�(��K(/�G�(��D(/�L�(��(�� ��~B��O�(��@P�����/��}����Q"|��B"ȼ�{~�J�*H.z&��F.���/t�����M})��H���j@/�j�/{� ���/�H�z&�/y�� >}?�}� ���Kx& �� ��32 @R/�����KdS"@����&���������!�U�
F.�!T �*H.

�!�k U ��F� bT��H
�
 � ��c��Fwњ�J>

�P(�<��ۃ�P@(��<�(�碨{�� �!��&��� �O��P������ ��/E�&��&� �� ���Fb�o�K�vˁ{�~v��uɨ���/t�� .s&z�? ba"⠛�!a.#�/�r�& "&!#&q�`.�.��GH"�ba�(/�H��!�&�H��b`�G���&��C2����J�I"�d�ƢI�&��p����� �s!rosr�l4��J�I"�dㄪ ���4!��`������B� �� �!�6@'r��H�&@�&n��Hbp�?sA�/��&���G"��n&���G"��j'm~�:�..�l!��������p����p �e�	��� )� �j�u0m/ k�p"�#jk  �����D�/�J� bH �!.!d��� ��lH�&P'� �&����i;)�f���/�&C(O�z����6~�Gi+��$ �3��R�
C��BQ'6$�4� 0e,�h���  �{h��b�h����H~ʒ{�� P(�A"P/0(X��#t�K    A  A AbAA     �   $Hz�c��

�
P�(��@�$� �g�P�	: ���0�
����끰��Q@ �fe3d�/�c��/j�gi������g��6|)�k�yiȜ�q��b��H�&wij�j�}�� �B�o�=�LM3M=3MM3K=3\a3n?�<C(/�P�d���I�&���b�b:� ���/��;�*
.

��I�bP(�<���K=&>�*?b� �W�/��Ȁ����� 0��? ��/�l�Ҩ/��/�g����/�Ө���$�&%�&Ӡ������&��&a�&�0�     ���-�b,�b���$(/�(�%)&&*&'+&�Ҳ���((/�$�)%&*&&+'&���~w��|&u��   $%f&1b'`bJb�i�F���y��t�J�X����0	�lj�kp)"#f�l�j�k�P�!��_ kHb_v^&9&ț&]�����4�(5�&������   o���ț&: H
�
�r�Tt�Kl,���� ��O����lY^&9&��d'��K� � . �� �|׀���� ��� �9&��4�c��F偬'Co6'�J���{�A��f� �	fo�����V2��Efe3��/cz�\bSbcGD����-�&�[鵞&-�,0�   �����r��v�0�	l	�l��'�/�-�0�$  ��/�Ѳ!-����-&a�&-�,0� ��,&�0�	l	j � kbcC(/�P�a �(�����OnZ���n�a>!(/����b�&�Z�Ҙ� � �I4D��Y�&�,�V~�|��<(r)r*r+r�|́� �\���́���� ��l���   �ͨ��Ɂ ρ��g �
����'��'��|������������!�Ã�� �!��&��� ������h��h��h��h�o�?��t��J��   ��4ば��@�^�|&�k�� �
 YS �������O �����3���8��^b�b�li�(/���,i�� �
�lI���cT@J
�cTJ
��d�43N(��7�+b�j��bc(c)c*c+jk+d܊�0	�li~r�ik�p"�#[id�h�&-�,0�   ��(����n�n�lii�� Y	 ����������Ъ����' ����(X��(/���(���(/������W�j������b	c��+(/��+|i�|�tq�5d�b�o�bl!l ���s�b��bk�he�2b�� �"(����/�ؾ�|�2�J&c�bbb�j!.�/�b�d����w����w�p�|��ڶ�g�Cq�T�*�\��@   e,�h��� �������������&���K�����|&��Pk'�	�(����n���   �
��'��ʁ����[ p������|�~�hly�~�_�{ ���<b(��TF��
&�&
.@��&7
7
7� �F.�G�b�c�� �k�p��&��������������8��9��8�s<��8��=��=��=��9�59�7<��9RSDTUDVWDXYDZ�D��D��D��D��D��D��D��D��D��D�E?WCGwKOwSWw � ��@փ@� 4֌@� 1֒@ Pց@��@F� ��@Ɓ@��@����@F�Z0��ff�t�f����3p�e�� �Dbclv��D�~��ז ��H
(���j����l� >��b�8p� ?��"�����'�J��!��⠀���'��� !>��vo�b �� �� /� /(��C�(���(/��(����R�)b�����J����#6�#+��B��z��(�2����"d!)b�]�\�&�����je�`��
�
�t�����`g�Sd���