����   � �(&7	238'?3736135<z $$ $$:$$:#$$:<.		z	-8-	-##     /8  	 ""  #  		         .#  ##	                                                                                                                                                                                                �o_���lH��VѴl��<���H�6��L �}���}xɦ%����i�&N�E���T�������hI����!Ѽv�Q���}'ǉ�f~�C�IU�zP=�+�/��}�Gш|3�m�پ��H��fʣ�|$8�\6�; �ɺ��(\�.'-��$�^�x�@�;�K�2����Kr�(�{�oC��:��                                                                                                                                                                                                   �	�@ �^F��� 0�^F��D  �^F�� P�^F�D�r \�5C�� P�vF�����2օL� ����4��F�����@F^�����@�^F�����@�^�����@F^V����@D�^���BB�^F\���@ �^F� ����� ����� ���� ���� ��������� ���������������������������������������������������������������� �  � ��N�ԱD��N�ԲD���D ���˄ ���D�������˄ ���D����C�����������C�����������8����5����� �8�eߋ�����5 ����4 �����M����� ���������TA��L�G�#�������������	����9��������7�����P ����@ ������@�FW���S��FG��8 ��FGΆ�8�N������ ����� ���� ���� ������,.(���� �       ���'��l��� �����6o��������/��������/��������������������P p���!�扮½�c��d��6��B��b��l�?��s�!�Ǩ?��� ���D������>"��j$Г�Q���$Փ�$��q2 ��i`bgid�i����g�J��J,�����iB;�*����@�� �q ��"����l6�m6��6�l�B&h6C��lʄ�Q��Ũ�$'l���x����-Y�$'����-��m�*-�-h�����/�()-K�(��+,��j�h�/�Ũ��� � �i*)-ś ����ʻ�C��#� ��8�L5`I�C � `B�T@`��X����� @o�� ݦS1Iw��0pm lR�H����·�.6sX�<��2b��i����ٍ���r�����Ȅ�$딦+),���  i�Li�,����B2h�cn�co�c�߸��
�s v�!9�F���̘�6�6��3 ^

d����6o̣� F� �� �|� �����c�o����|� �$w� '�s @b�h�y�)��p@on ln�D H����Y0��s
����"��y�A0��~��y�A0��&q .��b����Ӛ�E0pqbD�!p⨮�p>"4p&�?2 �c�op�  r� &pE ��bH
���& �0� 'p�&�X� ��� &p� �r>�&��J��Ā �� �s�� b� �q .if`g&�㸏E X
l ����n�op ��@��U  �    q  ��	&4�&��	�r>�& �J��&��&ߘ���	ǘ>"��d�ߨ>�&�	����>"��b!�⠲�4�&��J��D�q� ���	&��&��!	� ��>"��b!����4�&��J� �����b�@n?��׉�� �q .��b	4b� �                       ��?n�P�� �f�b���ccbG���6 6cE 4�& �̉l�� �(/��������������� ��/��cb��b  ��b�k�� ����= ��&�̲�Y����= ��&�̲EH
����k � ,�?(O�)_� Pb�i������Y �K()�E0H
�)-�� �.\�5[� bÅ?kF)f�� �a=�`K��  .˽�˩�����������˪��������������������ȾjcD.E�4�&b�bƽc�����cb��b  ��� �  Dbn�cb��c�h �O�쐴�c.�b�� ͸� �cD.E�4�&�-��-Ǡ �?��<e�4d� ���;�"�!i�F������;0H���o ���'�7�	�t��p��U uT�%�R	$)H�4m?uTRe�-,d ��>�mu�U�$S�R
 "�H�mu�WM$ҞR1*�R�mu�W%՞Rh��\g?3��WN#��Ofy?�I��q[c�݀�/pm?u����zm?uS�ME�$"/sͤA�p��/�z ���mu�W&�b	&.�f�寺 ����mu�Y�$Y�bf廵}�9P.y9�H��m? ZM�F�
" �/�y?�I��q[c�݀�/�m?u������g?3��WS#��/�m?uS�M�D�5"������mu�TM$�R4�)�1���mu�U�%��R+i6� ����y��I�Հ���	�;33C`3t�J��U��� n
�i����
b���h����
���|���g�JO`�gib;i&�P�z'��DNKw �sO������\O�$�p�}�9�R���/.gO3��WQ#��/8tOp@��B��P�� ��b�����f����b5�}�8\��j��zd�%�����qM�e��1�|v5�m�
���izf�}�8\��i��b�"��u����u���e��)�xx���z�fd�%�����t���}�X\�&�ܭo������� xs�e�� ���"��f��i�O� ���"`��/����D.��bH�����$����"����b�����+       ��!��?������&�&�&�&��?�/�.��bЊl�
�@ ���'���	  �/���/���/��?��          U
{�<���	�������	�� f�b�n��f���(���/���" ��(����/���嚀����"����H.&/���t���������&������"����?���h�����h׀���h�����)���9���� ����)ـ�� ��Kꀞ�+� ��]�=蛮��S �뿾�?���A�]�� ��/����/��b�c(��(��������︻����6��&��9   �
Cݤ�@����F����������D� �  !�(?�����D��� ���?��?�˻���W���b��"���@�(����i�=����c�/?�� ��QT ��� Jq���� �O�V�x �&�(���p.oN�� .�{���@�����P.�/��K�����&�&t����ǈ�(/���(���(/����Ǹ�����(���(������<�����&�����F���|�"(���kX#
�, ��#�� �.��qߧ�W� �`��� կ
F� ���6���"���¨�� � 
.

����� � (���� ��(� ��(�(�(�/�������� �����o��)��"����.��k��"����,�(/��������*!��&����&� ���c��F��É�ȁ�É�����뢨��� �   ��(��(뀸� ���}] Q��� ? �I� &�������6��)� �����)�������cb�����)�)�)� �	D�� �	L�� �	T��N7��7PR7 �4 �T��D �D 7      ���l�ˊ��(?�����������Ѻ�2 ���J��+ ���r��{         ,�}V�v�` �� U*q��!J����od Z �	�� � ��/�������ŀ�  ������ �	� �� ��6��'��)�&� ���4(����� ��b ����É�� .�/��� ���(���(/�����ǉ����  �����i����� �  �������  루��  ������  �	 �   7�/Dq������� � ��X̎3�K �	�����涃l� ����H���b��i��/������.����@N��,� �� n��&�����0��d��0J
�
.
�� �    ��C���P�`�V`V�`�Li!�`�`@��k�M� �������ҋ ��|���ỉ��ʀ��&����3���� � ��?��q�T ��'�����  `         ���� ����� ���c�� �� �����e �줈��  �¨������ �$H����+,��� ���ǉ����;���18   �q� ���&qD.
��
"t�
"@�����������$���������{ ��V1x̀�_�O���y�����-�<-�~ ;�� �b i-�� b�$�����qb ��i`bgidi�,�����i*)-��,�g�J��J��˃i�;�*M`�d��4�ʂ!���@n��"�����)� ā ����� �   ��'��'���6���b��y�c�b��{|�0 �      ���[� H0 �/���) ��Yo ǩ ���� ���    ����(���(/���Ё���|�6�����6�(������b�����!�������ÉΘ���F.������|�<�(��H�����!>��<����[���e���]���n�� b�$@����&��(����)��+ ���ǉ��a@ȿ0��:��U�[�8��3�P��  �] ���� � �(����bF�����b��&��É���� ��b��&�J.����b�ۖ����J.P����U����"��b��&؉<�@.�/�����&��É�Ơ�� ��b���� ��ے�����)�����; �         �?���� �         � �KNUk�U������P���� ���?�������FN���&��,��|��C����������i�����i��������(�����G �&��� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d������ ����� ���� � (����B���ǉ�� ��������9���������>���������ɀ 5���K(����� 5����� ���s!� ���)��)��F������< ������~�f�i�/��́���3���&��J�*���G �偼�|�Y��`�ˌF��:�?߇( �UN�<1��?  ��/�����b��b��g�'Ӝ'�����y�&�|���xE��r��'�>�����?�����FӨ?��0�����0��s(���tƠ?��������������� �	���(������<H����)��+ ��bg�J������|؞� �-�������0� ?@�-�v������k��ߗ��                                                                                                                                                                                                 �;��V�            ��  6�	$��2��"��$ �o���f��f,�t �D �v��f��frdJ'uIG�6�  4N   	    8 ?@ �� �� �� �� �  �J`HP`��������������   � �� �� �            ���   } � � �t 0������	�yr�k������$�����$��!�F���^$�����$ϑ!��F��b�$ؑ"��qnqD.q .tqb� ���s�����'��'��'��'�ʚ��'  � ��$���ʚ���w�$����ઠ����r��r߀���w� ��� ��� u  �P1Q���s���f�O� NRT���C�a���4��g.���W������]�.HQ�m~X.~�����i��(��f�<�Ƀ��Q�6���5&)cҌ�"bEz]�Y QT�Tay�K*�s��f5�"�5Y���c�Y�j�C�d�{�30� ��5h�SL�.��=�GR_$�؟tKRg =�ܟ��Q,�T��XZ
]! 	/�nvR��v                                                                                                                                                                                                �	���D6O>����z���/S���<�ę+��Vv=�o����Z�.
B&���l�� !eQfi�C�~��F��cm(c������\Q��X/S��R�5��~;z���;���I�pܔ���T1g��$
��ai���ޘ�)4�!���)�`�	�^�AM�3!�ԙ��%���_
��:^��)\�1��7                                                                                                                                                                                                	�E;�iثb/��A�,�à�-4��H�qi�!��-'�֢(D���FM�{�K��8���U��:G��(�PL�iB:<�P����%��?IP�)�[�,1�ݚ���@��<繦�"CHwX�E�n����s3�ԑ�����[�'.�\���@,U/x#^-u�N��={l�su@��                                                                                                                                                                                                .�����q��Ҕ�)�ƽ����S��U�^8b����%/v.%LL��� �~������L7�}X _�
/�OL('�%��}�W��`� ������`6��N���9'٥�'*�RI+q_l�#��c����Tyy��)v���=�7͐k�S��S�ڍ�D��M� �N{�����D]T���L܌�,$�B &�                                                                                                                                                                                                yFl���Ҥ5���F��8��Y<ɮ�v��>�2w��xf,�>|0��8k�ɘ�ggIz'j���_\�R`�$�����\;N��]33 x���T��R�=�|�s�7[�(ȧw^(4�($^�7���4ÂAܜ�1+�3���m9['��k��>{~�Q�Ra	;~�1[��>P/L�|8�&:����                                                                                                                                                                                                `���N�T�\DJ�#���tcծ�3����5`��+�6m'enl�SE	-3��<w��ۇ�U��?�pd����٣(0���G����X^l�-��'t2-GB�q�H����� R�I�����R@V$�IWZ"���Z7�1$x���;��]d����@�ǇfJ4�L�^U��pu�Z���Na�9����4�                                                                                                                                                                                                ����c?$t�,� �G�4�r|M���	��K�m�܋�ƚ ���>+�*�5$lP!���P���8b4Z�!"� N���B������C�T%�4"#�p��`1My�'g���l8�����Mh��d�B�0tXJ�OGN�1�Y��(ߟ���/�|�Z��VP��I�����ar�v��Y�S                                                                                                                                                                                                ��ES�k�*6��~�;nO���!
N���w=H�?�f��ifcL��.,�y^�6۾p�eւ>N���o�<Ǒq$��M���������&��#Y1�
�&��j̆.�{�@�nU��~S�y5��6�p\��L�B���������k#�x��2�� �Rju�%߻)o[X>,��!;�O�Uޓ������                                                                                                                                                                                                l�=�l�?�C�_�j�7�P�@U]0��)�_� UX�wk�<�o���
�	
�_�l �Y(_<��b��f&��'��t����	�_F��(�+hnH("Vt��Ox�0Qp�@@�F� K�f�f u�/�ԃ�;iC4�M��#��[��������
� ���Vmf�_��6*\*����J��ȓ�H�����%�                                                                                                                                                                                                   �b!����>=���& �
�������Ҫ����!�/������!>�/���������!�����6� >�?������c!����/�����!�����6� >�?�����!���� ���!���� ���n��&��'��'� �    ����������buj����9�( �	����b���Ҁ+ ���$
� �&��� ����a.Ӑ/��K ���6���� ���cѬh��K ��!.�H/�q�֐/��N� ��ʂιk ���&پ���K�΄�ص ��� �         ~ �	���ߡ� ���홅J���'������Hs�|���EGq�]e�ۨ�ջoϠA�Sjt�j �cLqWFs�=|Kr�h�
�Q�om?� �����2؅
~�K�z�RN1���A��lc�H�0��e6m��b��e��a����"�J-����G	:���	/��?�����#쀇���u��j&*v`�K��%�h2 9k�~+lꦙ�~���]CQ�u��ڣ��/ܰ�y/�����z�23͈o��kj2���,$� )>��0� o%$���*$� )0�;o� ������m&�j��nb��b��ɠi�
���a��i�������7�Қ����b�����(��t�������� ����d������j�&�
&���֪
�J��z��3!��� � � ��� Yl�+ �Љ��@���� �A?ݹ�D �  ��& o�
c�ט�9��b�ט�/�e����(���4"�Vnn/��s��y
�6
�<��n

&^&O��H ���������װ�o>"
jb��i= @�&(?����9�ܘ  ���J� ��
���� ��4��l��6��C��d������|܊���� 怼�� ��"��/�l���� �(�6�� ������V��o"��i0��'�zĄp��¨������h z�p��¨�u�����h z�p����il'l?"
jb

r:
&m
'm�+ (���pF��6$ ���K ��b+N�(-� s�� �۠�#Ӛ��jz6� ���6��)���   ��K 	��
�� ����\�� �����k�y�(ώ��4�&Vn���S�'��ő�� ���i��b��/��� ����/���YH/��������龽b��&��"��bF�����b����D� �       UpHb�p�ƀ���k ���(�y�� ���b

�
X������bF�	��&� ��Pnl�(Y�lc@��lD�
�遬������������"�������c��c���	 D B �AD0RD  �P ��'��'$՞����q������'��'��0Q�'��'�$���阶���$��������'��7��'�$�����7��7��7��@�b� 0�# U �� �MA���5����5BR1 �BR �;�6� �������̉�T�����@xD�	��,��@��g�n,���3�L�wN�S%�&�ul$q(.^c%�#����gLX �𡉅-'��
� n�vƪ
�.wD�$�B�t������� �|3-���`6GW����r=׭��2��t��;��p �]$��S���u_�J_���}?+�N�G�a`#}뒛�o"��,�0$7                                                                                                                                                                                                ��|xc|$%�d��3@��=ʼ��暶�ɨ����̌�<(��P�IN^��H�;B���;�$��r��$=،��E�Y�b@�������~����~�gn��-"^�7mM��l��}
h��I�C�1�VC��!�k��#B�l?ԟ'�kGO'�W'��T���:X���i�x�O�j���DP�+ �����                                                                                                                                                                                                