����    @� ?    :    ?     :     :    :   ?  %## ? %##-8      :   ?  %# >    ?                                                                                                                                                                                                                                                                                                                       �7��@� ���Ѝ��ưt�W��?�������F��� �? �i����!�l"���  �C�5 ��8���@ P�8 � �� .� ��B:D)3D#�B-�+i�*�x&xw)'�/��+)"vi  vI  
vI  
��*!.bw��v�� �u��|��*D�{����*�x&+)"ti��v � �v � �v � ��*b!�w)'�/v�� t�v � v � $v � �.ui |	�*��J{��� ��)�s�)br�&`(� `t���� �, ��.'f�q�p�)obnb)b�s��n+)"bw'��v�� �w)��v�� u	�|�'�D�{���� ��!&��&��&�Ө���-��Cm��(��Ү6�-�-�������������?�l�k�j�&i �}�m ��|���/����l�h�&i �}�m ���0���|����K ���. n%�ol��g��j�f� �bg&�Jz	�q)�q�(��!)���p)&z�B�be�/�ol����f,�z�f,�f�!,���z�)�/��(��@d���!.b),")b���z�c(&bY��_w)z��v�� �w��v�� �u��|��b�YT����J{�������� ��/�l��a��+��f� +����- N`-�aY��K ������K#$f)D._���s�`y(�`&��`I!�`��`I�`��`I�`��`I�`��`I�`��C^]"� `�ai ��d\&[&�O��D�O���ai �
gqD}�D��D��D��D��D�<B�i;)��D�� ��Zbb
�Y�X�b�Y��W �(?��V0'�JGIJLB6�  ;N   �l��f+��ޫ&&c(&%)f0.f�n'�n/b(���"&U�� ��6�@?��T�&)r"��b��d�6�B`n(& `B�/   �| N�J). �d�!.(��b ���ʫ f0�n�!&bY��_b�Y�O)r"��b��c�d (�%b���'B.�z�A�! ��<��� N�J). �d�!.(���b ������㪠0�%�/�A��'�B��*�!.b)br�& ��b�Y�Oi�}��b�YT��   `"�aY�[ �
��)��&�@���E��� 0�H> ���6��d�>������� �S���/���(�������K��b(����/���� ���/�R������"���Q�*��"H��P�*      ������@  �o/���&!��"�$b���#�J��O�/�#�#N"����$�M#&�R�&!��L�&!����#$f� ��
6��C�d�6�
Ct��(��H��� ���6��C��d��!B�螠B �ᒀ� ��.���� ��'� �   ���0 �������� ��W��F�響�� ��D������K �F�Ⱥ���K ���"�����&�D.���b��7�.��4 ����+ecM]cM��aG����~� c	���TR���H�c��҃ �N UR���H�c��T�`R��D��� �� �AA ?   R�z f?   Ԅ��40� � SR� �f?   ̀� �f?   ��:! �?`  ��@ �?`  �� �?`  �0 �?`  ��� �f?   � Q� �f ā: f ��: f?  cϘ��/cҘ�x+`�S� �S �S� �?` c	CP`� ?`                                        X5��q"��no�#���]��s�ir��r3�&��Sl�/���� .��b2�$��������//�,C�X5 9"),F��������� ��WWb� ���� �[[b���]�      [�   ����3 v������
�T􀓶LT&�p�
�b� �&!̕"���� /	,C�X5 ��b9"),)���t�&��vK�&�)�����D�/�/,�C,y1� �!^�U�n]	&v�/�L�T�np
&e8 I�&��+ XX�-�������bO�bPOcQQc��QOtP�J��������D��Bp5jcU�SM,6"%&!!.�Z����rb� `��<��t��   �MN ��A�RA��� 0	����DG�S%�RA��D	�T�`R��D�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C V`!ϔ� C�TS���@P3 P̀�D��C�À^�T@SXGS�TR���@                                                                                                                                                                                                