����  @ /("$: : : : : : : : : : :  :   	   	   	  	  	    	    	                                                                                                                                                                                                 
           @�   �ܹ� �D�  �7�˝1�'������ �@��h�[U�GO�`��d��ɶ̞��ih�P@�h �   �  F  � ���?�U�Z �� ��         � �                                  �	'   ��
�Ĭ��o g���D�������mmb��&��,;�r<r=QvPRfS `�>�:�o�:9&XWfb�n,؞bb9))%#����b,i%�� !���
9")(��(��,�( �!��9")��"Ӛ,��"����9))�"� !�� WI��
 !�� �g�6)��
 !�� �g�6)��
��� �!萀��  (?�����Aè��îg6b�� �! ��[�\[bg\b#��\����[[b���\x"��� !��6K"[�n\\bg[b>���[[&�[⠩�\�/�\�� �!$���l�v�&A9"m))+)(ʚ�@�b%i#���,��b�%#����g")(��خb%i#���,�b%i# �!?��                         M[&\��]i^n_�G�Fn&]g&\)��_g&^)��n�J[�J !�� W�o��:�����:"����,�ob&�:"[�n:\&\")%�#���,�\[D� �!�����,��:[&�:�\<bob&\"A))+%�#���,�ob&%#�����,�b%i���\[D� �!ɑ�� .�(0�:D�L����� �W6B
[&�,��<�b�nA9")[�+��%�#�����,g�))���b�%#����9))b%i#���[�� �!� ��!�	Jg&A���giA�* !�4�*E[&H)Jg&[K 49r54sb���g&[K b��H����[�� �!D��䫀S"�}�bjdb!.�?�r����=��!�z�<"�i;)�f�Zm�E[&I)Bg&[K 49r54s�����g�[K ���I����[�� �!���E�[Hb��[K 49r5Jrg4c���[�� �!����E[&g&[K ʒ�H����[�� �!���E�[Ib��[K 49r5Brg4c���[�� �!˒��E[&�g�[K ���I����[�� �!��E�[HbÞ95'�J�g[bK644s�����g[bK6��H����[�� �!�������>,W�NX&YNbTSf�$��P��g�A�Y�| T�i P� Q�giA�:��) !�/ 0�,�WNbXYf S�NT&P�i��g�p�Y�| T�i$���g�P� Q�p���Pgfp���� �!J� �τTՃ�8��C ��ix_�bE[&I)�9�5�~Bg&[K 64'49��:Þg[bK6���I����[�� �!���E�[Ib��[K 64'�9�5�~Jg&49��:[�J !���:E�[�ng&[K 6)��:I)���[�J !���:E[&H)�[�K64�~95'�B�g4c��[�� �!ԓ��E[&�g�[K 6)�JH)���[�J !���:M�[JbgLb%��,�v�&g))8*)[L +\�%B����\�J(�����[�J !��JM�[bgLbH��,�v�&g))8*)[L +\�%B����\�J(���[�� �!&��E�[�n,�Jg&8*)[K o���g8b*[�K	o�Jw�&�,�abf-$����[�J !�K�L� 3	0��T1)0 �U1)�=�khwE[&�,�H)Jg&8*)[K ����g8b*[�K	��Jw�&�,�pa&qb&-$����[�J !���LE[&I)�9�5�~[K 64'�J�g4c�[�� �!���E�[Ib��[K 49r5Jrg4cؔ�[�� �!Ô�E�[HbÞ95'�[�K74�~Jg&49��J[�J !���J� � ��� ��UUb�_�E[&H)�[�K
49r5Jrg4c��[�� �! ���E[&��g[bK6,��I����[�� �!���E[&g&[K @��I����[�� �!-���E[&��g[bK7V��H����[�� �!A���E[&g&[K 
)k�ZH)���[�J !�W�ZE[&H)�[�K495'Bg&49��Z[�J !�l�ZE[&H)�9�5�~[K 64'�B�g4c���[�� �!���E�[Ib��[K 
4'95'Bg&49��Z[�J !���ZE[&I)�9�5�~[K 74'�B�g4cʕ�[�� �!����E[&�g�[K ޕ�H����[�� �!˕�E�[i�g�[K 6)��ZH)���[�J !���Z� �y��ny��{�z��E�[�ng[bK
��I����[�� �! ���E[&�g�[K 7))�jI)���[�J !��jH)49r59rmJ"g8bi�nb4ch8b�g��4���ݿ�eebB�/����4�у�gg&�5�55s��4�x�/� �!*��ޫ� `{&T&�7�O�ߣ ��J�B��/�ߣ�z?'��K��@	�0T� �y�[�m"9g&�/�zf8i&�b�[h&8�-g�-[�-���e�eB"���e	 ���v�&�y�����u��Hb���[����gg&g ���[x"��� !���j�y�[\f9"mg&8*)g))[+)(К%B����[�J�g�g\d\�/�[�x�/��H)�u�v��o !���j� ��h6-���C��ă  �y�[\f9m"g8b*g�)[�+(��%�B�/�[����gg&\\B���[x"����H���u/v�&� �! ��D�_i]n^�^g&])C�zH)���_�J !�4 pD_&[��\i]n^�H)^9"5]r4\rg[by��^�Bg&])y�z\g&[)y�z^g&])y�zH)���_�J !�P�z���F_&[��\Hb\�95'[4'���\�Bg&[)��z���\�g[b���H����_�� �!����y[f\9bmg&8*)g))[+)(��%B����[�J�g�g\d\�/�[�x�/�ЪH)�u�v�ӈo !���z� � b��'{j&Tr&{&jbB!���b .brd�T�(/�!�r�kn���/��r��ޜe"Zm�7~�
[&�_&�^�[]&H�*^H.�M�
["]IbE�\`f`K 4]rDE�447��95'5B2g4ce��`�=`&\�J^�J�c��^�[]&�^�H��M
"[]&E\&`]bDE�d�og�`K d)e�c�/HH"���`��`&\�Jc^d�[�	[&_�J !�  ���n �T&{&N&t ������}'�J� �  �,�P�WYfSNbX�nQYb| T�i$���g������gi�����) !�� �Q�k���:(/�!�9�/�Ԯ99&������93i0W��,�WXfRQfP�k��>9FX&WHb9�54wJg&���J�gi� ��
�bvb�eb#�����,�g&��H� �!Ԙ �4� ��         ���i_� B_:b ^�]]b9]b�,]�^�J]:b ^�])����]�]^"�����^_d�]�: .^]b�����]^D� �!���� C_:b ^�]]b9]b�\6\�?�\����0�/6),]�^�J]:b ^�])�ߪ�]�^]"�����^_d�]�: .^]b皈��]^D� �!5����� xLV2m�ح���:�� �_:b ^�]]b9]b�,]�^�J]:b ^�])���v�&�]�]^"����ۢ]�&�\6�	"�]b9Ibړ95'\4'5B2g4cؙ���g6\)�֚I)���])_��]�: .^]b͚���]^D� �!����� o )	g")ڞb%i(��b�%B������KC�/�ܫ�	�����|�|�T���_����[�nW8b8�l[[&[> 9o�\���]o])�[�DC���^[bDJ���[g&\)?���[�>5[g&\4'^�/\�?��^����]) !������>9�X�WHb9�54wJg&t��@�9))+%����I)Jg&t� ��
b&v�&e#)����,�g&t��H� �!Q� ������2;���ǯ ������Ȋ��)��;��6��N��&33�R�/�0�r�:�>0�&�60 �30���ހ1)�D>���0i�����a2)b1)����D.���0i�c�2d�1����b��b�b��b@��D����$��F0 �19��JQ�/�����������+��+���D����D�J� � ��d�   �ZCr�O� (M�&����ć�������(�� �llb!b⠑�� ��a�K!c�/�d�!b⠙�� ��M⑙f��J��J� ��M⑙f(�������������K ��eeb� �jjbijb��� �hhb��� �ggb��� �����K ��� ��� �VZ&�.�.���.Z����
.)hhb�Ƕ!?� � �.
�.f�fk&k�+ �VZ&�.�.���.Z����
.)ggb� ��8�Nbrgr�J� �s�n8&Or&s's .rt�?��{քo
�������,g��)	�,� �g")� g��g�,���   �	����%I/��*ڞ.-�'&�3��,O�� ��n9�)g�Am")ג+(��뫈���v�z  �P�/�T�~��y�cz�dg� m9")8�*��+��خb%iB�/�u��zG�t��e�	Q�/A�����g�DC���y�jv�*   b8bjgb�!j�?�g���
jjC!h���h�*�N�rjdj!>b�/�b� b�r�Jj?B!j���?�*�b�y�/��yvbz�~bjck�d� ��N ��`1��	�G@ �VZ&�.�.�.�Z�J�
�.d�VZ&�.�.�Z�J�
�.K�c�k ZZ.
>�)Z> �)� ���������� ��  ����&�> �)�.�枼J�)� ����ɶF�F0(��@�
�

���G(��@��)��N����@�� p&!��"����DM�P��HG1L*�����D� ���6��B�9bm))�,� �c��dg m9"A))�+)���b�%���e�@(/�@����,�g))��%B����g� )b�%���������t��v�� �  ���"��&�2��"�c��"��&�/�x������*�0.��b��&��'�	"�n���>H��� �o�� @   �P����� D ����?�������;Y N��6W�/�X����,����K ������b��b��c  c�� �t��J������\a�RL�AX�e?�H>f:Af<�f��f��f��nQTfW�P�nR�n,؞m9")8�*+����(��%�B�/ !�Ϡ�QPfS�k������������������D������  �� �TSG�S%�RA��D�MN ��A�RA��� 0	����DG�S%�RA��D	�T�`R��D�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C V`!ϔ� C�TS���@P3 P̀�D��C�À^�T@SXGS�TR���@                                                                                                                                                                                                