����  @=
6.=: =+: 
7,= +#	=+#+? =6  =>(/22/2e= =-&=f   :     8
8
8
" " *  <(. 
<(*
=
	$.$.?    $. 988,$. 
, .    
 8
8
8
$
 $$.,  
<$.70 6.:  ; 5<(/= 888
8
8
'43<(/2= 10'4+    ; '?+(8 //C/<    ??? = ?!  
 D   ?'>*?. 0==<-
/..<(*;>(*#-.*:> * ;'98'9'7 .  ;. ;6 
 �� M��� ���L �    � =	��	�����7�*��r�  �  !�@                          �� 0                  � 0   ��������   (0 8? �� �� 0��" D��D��D ����s�
��� �v���? ���?���R��` �������>���_�&������8?f�;�f�'� �XA Q�B�iB�/���!A���8�b�Br9I&I��Br!:�IIk�B������'B9"IIk��'�:�IIk��'�:�IIk��'B!.HI&I�@�"@�i��'@Q 9I&I ��!��� 
.

������  �`��P�����W��3��%��S��3��7���8�/����ں �<Mb=Df(�(RD&)�(SD&*�(TD&+�(UD&,�(VD&-�(WD&.�(XD&/�(=�K<�/�8�� ����=O���C�i<�K�C��&Ic���I�JID.D���� '����!�� �&��ͺ��� '����!�� �&�����ۺ� 0            ������'P�W4j B�?6 ��C�/�/�X�DJf����J��7���.�/�W�DJf����J��6���-�/�V�DJf����J��5���,�/�U�DJf����J��4���+�/�T�DJf�ʚ�J��3���*�/�S�DJf�ؚ�J��2���)�/�R�DJf���J��1���(�/�D�J�i���J�/0�K�?�?`��؇����#���������C�7�/�X�D�i�������6�/�W�D�i�������5�/�V�D�i�������4�/�U�D�i�������3�/�T�D�i�������2�/�S�D�i�������1�/�R�D�i�������0�/�D������ '����!�� �&�������=��!�z�� ����Z1��1,�e 	 ��D_"��b��s��s�Jv>.���>
.���>.���>.��� &������Kf�&!������B`�c@�� � �C#B�S�   ?�l??'?�J?!.?�?�?��C�_�&���?F&?E6C_"Ձl�D�_�&����/�פ�ף  kq�s)p&(?���A�o �4i)3�&����@L#3 N3%3 ?�?� ?�?�J?.?�?�?��C�_�&���? .F?cECb_�&���D_"��l� �?�l?L"??b??r���?L"??b!?㠾�?�/�C�_�&���?F&?E6C_"Łl�D�_�&��� ?�?�L?&? .??r���?L"??b?���?�/�C�_�&���? .F?cECb_�&���D_"��l�@���E���/5!�T���f�b����f&�����fn����f&Z�뀝�fXn�@�@@w  ��� C!D⠠�� � %����� ��J�G_bC�&_D"��b��bD�&�GÁG�G�<!G���G�JJ�/��� )*+D,-D./D�.�-,D+*D)(D� �/.f-,f+*f)(f� �� �AJ.!���� ��w)  J
�
��(��H�=�P ���6��C��dY .�J

�Y�!��� ��F.��� ֠'� �    ��/�����{���c��bJ
�
�跸(� � Y (�P /�Z��O�@����*N /�[��M� ��\/�)�����0 ��`c��C�`CN(LC Q�L ��/�`���3 ��}FE�d�8N���ヌ �  $�����/�Z��� �#����
�Q^��bLK&aK��B���`c�      �  	"��!��������� �&���� J�����c�re �r� y$�� �#�d;���b �JOԀ��c'�e' ���'��B()*'��:��i��ޔ� UG�S%�RA��D�H�@|� �������Ӹ�q_HL� FP�TR��RA��D�D ��0	�S  �JO����c'�e' ���'� �JO����c'�e' ���'� �JO����c'�e'b� ���`c�H� 8�� H�� �� S �-�k") �G� 諀�Y�����b}�k��� @7rF�,� ��G��ħ�� ���`c��x�E�hM��T��� ���`c��E �D&��%5�!���� ��/�`�c��L��T0O�#���N�� �F����`i �;�k ���`c��CL� �4�0 P�;�� ��@��ɑ�ə�ɡ�ɩ�ɱ�ɹ�����+B�($��+����+���+��� � �� ��_Lb��s����@���   �/�`�c �@.`����N(	�$��DM � �]��� �(0&)1&*2&+3&,4&-5&.6&/7&� ��/�`�cԔC�L���� H/�/����.������(-�/����,������(+�/����*������()�/����(������(����� �� �� �� ����'��:  	�o ����&��'��>�!.��/������ �   -p��.�" ����o�J��s?b-n��"� ���q����� ��+?�(��kabn$is^bo�n?-)o�J. ����n�Jan&^o&�?�-o��.� ���n������ Kr� Ғ��  0��6��'��'��K u !��&��<�rq�DJ.^�ai?aF�ayE�/�`�          �   dDJ.^�aiG3�/�`��C�� � `	      �;�d��Q�K����Q ��?/�F���E/���J
�
Q���d��Q�K����Q ��G/�d�V()l)))>�-.� �X����+$�kH.���ssbZkr)��)��!Ɍ������'�����j�/���Q�i�������'��'��'��'��'��'��'��'�� ��'�� ��'�� ��'�� ��'��'��7��7��7��7�/�߳f�b>l���́l�Z�{{b ������+$�ks&���À_353��#���d"o\!gN��YL  Z��� !�� �W���� ��┓b��d��������&������� �    �����&��⁺�� ����
Q(����/�����/ ��b���k� ����� ��b���/є���/�����b��/����b���&� ������&�&�	&�Á	� .����Ӹ� @� ���x��x��0 �8�? ���P@�܀�n����&�&�	&�
&�&�� (�?	�<Q�
ǎ����� ��/�� ��!��i ����b�i�v��s��}��m�� �l�����&�ڦF.���d���!�⨧�i� ���    �!�����}��y��m�� ���l܋p��܋����ܛ   �ǘ�����   � ���� ����Dh�����K ��
.�)� ��!i����&,�!�"�� � �\)� .�[b�����   ;�� �  ��������&��"(��N�/��շ���/շ����(O�@�淢�����c��b�����J����@/�R�H�����v �����-�'��� �m�� ���6��C

�
�蠎8��J Y (���(/���H��])���ݿ@  	�F��i�����K ��
.

����� �Q����  ������/��Ƚ� ����(���(/��������s . )i}C"D()>-)� �{{b �ҙ�� ���+��hi��ZK) �������� +	ks&s)s . )i}F"D()>-)� �{{b � ����+l�ssbs�  �)}�FC"D()>-)� �{{b �����+l�q[bpqb��qq&p�Jls&[p&}())>�-�� {&{ )����s�spd��3����+$��)�lZ'}F"(>�-��}()>-)�z� l�s b{ b �Y����~�/���)�h() �bO !d⠌�e!.c�/��K�}�U�
\&�`&�_�\^&K�*_H.�R�
\"^LbH�]afaO 3^rDH�337��:4'4E2h3c���a�=a&]�J_�J�d��_�\^&�_�H��R
"\^&H]&a^bDH�e�oh�aO e)��zd�/KK"���a�?a&]�Jd_d�\�	\&`�J �� p�2�n �      