����C� C   	 	      	  	 	 	 	    	   
     
 
       	  -                                                                                                                                                                                                 ��b��b��b��f�(?����&��&(?�������k��R����(�!.��/�����/����� ���    ���x��h���b���t�.��α'��D��̴�4�K �(��@���/�&��"߂l��� �����&��&�&�X��J��� ��唀��� 0����Ӆo�K��2c����� �7�
���`�������&�6��9�|��0�c�b����(?�!.b�c�� ��&��������bd�?���r&�'�" n&��0���!>�?�����������������1 � �
0` �`2����� ��݄w��w����&
c�����	f/�"b�&�&
�/�����(���(/���!������/���	����&	�/��#���� ����D����"H��� �&���!.c�������s!�e�ɫG�J��&� �C�{a���	a>���_?��Q���  ��È
��8@������������?�����0��a�o���h��J�&�,����"����)�J���!.����������� ��>������h��0���� �����b�bD���b����)�J�˛ ���ށL!>���ޯ��������������& gJ�pIQ�������"&6������������������F� �� ������!.�������� ��&������ ��[�6��r؉��ǘ�)������		c�&����i �	ԁ�	�9�	���� �� ��(���,ښ�a�9&�fI�̿�̂`� Jw�gXB��>��o��  A���B�����д����O��B��d� ���fҠ/����b!���	�����0�����β  ������J��b�$`��(�� ���b!��� .��f��B!����&��&���         ��i
�   �زӌ�   ��� ���� � ������d��6N��\����【 T �g�J`x �(���c�����i�/��
���(��d�������0J
��(��&�������)�ø���)���Ø��/�D���&� ������� �D.��� ��c!���&��f�(/�@�/����J���ԽD ���J��) ���Қ��b!H�ǒ&���g/���B
��d� I�� ��"b	�j	
&"��&�?���h&�?������਩���(q>�8���hq>�8D�J
$��	d���� �������ň� �!.ccrtD�ū "b&� �!� �f	&2	c!�����)	�?���&�ή I��OE	  ���(��b�����(������Ѫ(� ���{ ��,!�������(��"����������K &!�����  ��N�b�c���(�B������ !��h��J� � ������� �D����?��� �

�
�� ��)�)� ��&��8(O�ɨ��籸?� �� @� ��	����� 	��G ��K �� ���;���� ��Sem >L#� �L��1 �:P��_  ��SEm; �`A���  S�`S ���OB�Q1AS�O�#� � N$ 	Q��@�@6R���ETN"�� 0R���@�N2�� 0�8�`3���5TXL@!R���DDN�N E	���@a��PŃ��C R�XRC!�T �  ���1�A�P@�AC@�b��2 U0�� �C �S�Q�R`S(�2TK�$	���8XNR	�O6RXSe@ 0������<�������c�߆�8a���ؒ�c�a�0�ś ����0a�����"���hY����F ����������֮��������P�����(?��'�&��)�(/�������J�&�&�)��/�֮ /�/B�����������"����b��c(��������*��iT ��̢��r�b��c��� ��آ������������I����������C� �������Q��	���1����