����    @58>4(v A 0+ 
?% )$"1? 5?80  #!#$   ?3, 88 = >
< ,*,0/9'>.?9> * )2>2? ?  
   �B B 1���������                                                                                                                                                                                                                            �+&@ٔ�MA    ���                        �                        ��7��@� ���Ѝ��0 ���� ��dǧ�X�B�� � �XU�υ��   ���8� `��J *��˹g�.����j�P�r
�� ?�  
 D B�FF���)�~�}&���|��{iz);ٷ{A���� �yx� ���<w.� ��F���h�+ ��v������� u w$� ����k t	�Ê�Ϩ���� ��@.�/��B� ��@.�/��B�s�� E���`TpBR�� s	��TO�#s� 0wu�|)�ظ� �� ���P���?�֣��������X0��� 0 �/r~��w�r ��
>

�����q���K v (��pv p&w,�(/������)�o���n�m �o���q��"淑���;T�B� w����B3R�8G  y����� 5`���PŃ��I	�� @y���o��R1��D�8S�nyC�rR� 8   �� �}� *��*�h� �lk)j��� �i��kj���� ij���	�i��kj����	i��� t	���*�/xh��&��&t���Ĥ�s��N�TA" �0MN0 ��0�y   ��&j��� �i*������'j��� �i*����j���	�i���	&�
&��&	
7��Jj���	�i���� �� �  ���?�����d��yށ �gs�`��`6NR�NAD�E3��`Q�`VX(�4�T��C�s�`�N0RM�`P��E8�8I, s	�N�Ճ��H`2l0� ���`@� �8ƅ1�s��(�U3�� `�S� NA��Ec��;s��	�#�B�XC�`�T��T0D�`��DE,! s	�� U`�8Y	N���R	 sYS(T "`� PT5R�RA҃b�;� ��f��� $e�&*�/��"�{ �	f����e�c��e�B��&*�/Ȼ��{��: �	/�&�d)x��c@./�/b/��/&��� �i����a���+�/�t��x�/'��&��� �iʻJ]�b.�� �� S `	������h�� otI_�/�h�O�����x ��c�(O�������J�6����s��� 1��TO�#�8�  y ���(� ���&�(���/�f� � ����&^0}�/��t^0��/��]���"t�'f@�@�����b]���"�{ �8 `������ ����  � "}& \iz��qO�}O1v�sO�O�O�eO�kO��O�mO� @b��/���t�o���q��)��^(/�[�.b���Z).�/�Y��.����X)\z���r��}1� .�/�Z����^(/�[��j.�/�Z�q��W� �qy��[&qV��(U�󚥡�%�,��� �+�ht�T���&+b^�b�F�D�b��j�h�+ /b� �S��S����"��b����D.X�泊l
�    R� /ʲ���b��f��     R²�b�j�bb�&��b
�v���$$b%&%�<%%b��� ��&�k ���d���� ������ � ��P� �	(z)���������������       Q� ��f��@ e�&*�/��"vt���*��x�P(���D.F.+b���O ���f��?�e��b!����!.��y�s���� �`1��SE`�	E� 0y ��n+ti�@.X/��+b^�b�F�&ီh��H�g�}Up� ��*� *�x�t���P�(��+b�x�N ����M)�����i�� i��&�H?����b��y��� i�s���� �N3Ճ� 0y��s����S���OB��3̀ y �nȖ"�/�Ӳ&!�π�� ��  �s���.�H�8Մ3 y j	��7i��2�����)j���7�i�F>w�7f9�����T�� ���ň   �t����*�/xP�(��+b���f��?�e��b!�4�y��!�����K��8L.�$N��O��R�� >m����.o����  ݈�B�-�$��Ҡ��6�����=m����ѝ�o����� ����Rc�i�󇭀 � � �� ��   �4�#��g�}Up�u �	��	i��(����	�i����+i��(����+�i*���.�l��(��ɀ� i��(���� �i�� ���0b��/�*��w��'� � ��(?�ж�*B�����7*�/��D� � � ��@� @��)�մ��&j��� �i߲��c���� �j��� �i� �Dbjl��BQ�)�@�������o *�x�a(�x-�-L �b�g��,�hK!��hK!�b!�(�����&�,&����/�-�F�,c�,�z ,,�"���,^0{�/�,�
�v�H(����$�s�`ГRTO�#� 5E eM$MN Qy|�(Jitz�F �` �S?� xs��� G"(�@�D y g	I������`�����|�t(�x�����h���/�ݦ��bc`���/����*�6�6�c#*f)&S�����)&#(?�#�d�##6����#���/�y���B�`�H(�((/HG�(|i����s��N�Rנ3TBT%`��A��P  �   y �*�N|�)�k�����*#)B�j ��#&� �   &ƙ�q��S� &(���ji�� i%u �&(�/��''c@F☝�'(?�(����'�*s���� `[��	��D�A� 0y��s���� `[��45N�R y ��ji��� i�s���� `[N�Rנ3��TO�#�8	�$�#�4y �@VO���DE�� DJ��Ān�� 5�T@0�                        9 �?��B���;��7�       �	��ɪkɱ �      bB�kY�qM�z>��N��ʣ          � �� ��  � �  �� �ň � �� �  �� ���Ĉ� ��� ��  � �� �  �� �  �� ���Ɉ�Έ � �� �� � �� ���̈� ��� ���ψ� ��� ���و � �� �Ɉ�و � �� �  �� ��  � �� �  ���Έ � �Ĉ � �� ��  � ��  � �� ��  � �� �� �  �� �� �  �����             � �� �Ĉ� ��� ���Έ � �� �  �� ��  � �� �  �� �  �� ��  ? �F�W� �	�� �� ���?�(�z������� �      Q��s���� FP����LX� y %Ȫ�s���� `[� 5�.N�R y *�x�`�b�����'� ���FD�*.��|� ���DD�*.��ˀs���� ��OB�3RQ y E�D���F��F` ���� �	*F.����{ �	*F.�!�� �g*������'� ��f��@ (e��&*�/��"�{ g	t(�����t��/x��*�/�"�f��@ e�n&�"*b����"b���r�{�"c�r�{s��L#� �Q y+�� �� �  ��O����? �,� 2�Q�� ��^ h����
 g	f��@�e��*bD��&7�s���� 5`U��HA�M�`��Ճ4@y g	I�� ���4(��!�`��D.����h�!.���� �{��|��� �             9	�G��Ly�Ty�?��Y��^���� ���������9&����Y��i �y �f��6� 0            ��p� �f���� e��*b����'� ��f��� �e�&@>w�/e*��Y��'� ��I�� ��׈C �B�m"�B�f����e�cu�b�!.s�{ *�x��P�(��+b�x�c �b�� ��(�z��������������� �      Q׻ t	��/젾|�    C*ڪ���� � ���&��(�.�攄J� ��CA��      ��4�&��4!!�!>�d2���!�J����+ *�x�a/�+�/xt�b(��� /��/x�� �%�/mm"@/�b�/�"/b���a�+�/�t��x�/'� �/�8�)~�6~}��b~�{s��� 1���yRU��A@�(D��C�� *�x���)�bd��)��bdx���"��{ (z�������������ϩ�ϩ �      Q�� �*�/xI�� ��*�!���{s��N�Rנ3��ă@y *�x��P��(/������� ���� ��� ���d��6��C(����&��7��D� �    ��uw�#�:�8������� ���DE FL MN TU VW \] ^  �hBL�D���a����/>���bń��'��'}'�P � ���(����@�  �i����b��y@ � i� � �����   �Ȳ��K *�x�a(�x-�-L ���-�"�b�-F.-��,&�Λ��/�,��-,�zGĜ       R�	A����J�(�                                                                                                                                                                                                