����     A: 
./
 ./1!  8>(*+?7<: 7:8 
0>(*);7<: 7>? .:
../
-./
?  
7"9
8"9.1
  0&0!*;: .9  0+ 0>0&0!+=<(/<;<(/:9<(?87.?  ?7>(/65/U5 ? 2>>?=? 8                                                                                                                                                                                                ���v&xş��C ���G �   �� �� ������E�?D0   �&���(ˁp�   ���8 �t�C ���0���7�@  �   �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s�
��� �v���؇?���������ȶ�@�JA�J���!B���&�(?�B�����Ĵ�6��C��d�!>C�c��t�CD�����6��/@�����"��j      ��2�����2�����&��C(���������C�F�۵d��0��&��C����b� ��!��� 
.

������ z (��~z ~�/?��� �yW� �S�_oQl�l��	 �Q���  	��A���� �Oj��jd v�O"�p
�
��� H  �y |���D�PQU��A	 S ���D" ��P ��T                           ����������'��'��-������ڭ���������  �  ���������(��������t�ګ �B�������������K����?� a� � ��݀������ٸ�!���0��O�٨����J�ъ���ǀ������@  ���J�
>

�堮��c��@��b���� /��@� � ? ?`��؇��� � ������� N�������� �H/��O�������j8�   ���ƌ�+	������!����̯�&�����"��hˍ���&��&�톖����ގ���"��* ���O� ��F.���+��   	���F�H��	�������j �
'�	a� �����᠎��&��(���������္���� ������	��F
�������h�� ̅ � ��� ��)��)��)������y�zzr{�}��݂�چ����"���Äڴ�툉���r�������>���D����߯o�1&"01�1����++���,�(�1�-1& 0&�+(d' ����+�%� }�9���N��ߎ��ڨߑ���ߓ����+��B���a������-��� �⨩�����������⯭����P� �(��(����  &!̻��� �����&!����(���(/���(���� � ���-�����'���� �M�/|��� ���y����J���� ��|�����A�?r ��_���8 ��)��)�����������F����������y�����������(��
�����ڎ�҇����� ����������0���?�I�''�'}������~ /�ӂ�*���
� �    <aR��b��&�K"F�H���&�P.��/�󩀀�S�����G��P���� �?�1�� 9�P