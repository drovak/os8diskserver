����  @ @�      %1.$  %1%2 	   /  %1%2   %1%2       /  %2..  /(  %1%2  /.  %1%2	   /5x   %1%2                                                                                                                                                                                                 
 @ٔ�MA�� ���L �                                                                                   0@ � ��  #������ ���6�W��$BV 2� "b9"�)"),A �m� t�R����"��"��?�R��` P�xm���f!��/�,�������n)�n)��(����n,�F .'Pn'�'�' !D�'"�jm͝ �o?��qif!��/�,������,!.�(/������n)��� (/�Ы��,H 
�
�pf������,F pif����/�,��Gpi� ��� �� �� P �(?�r�� ,
D"�bnȒnȒnP�nf������,.L�&pf������,D W�/�,��Q�&pf������,D W�/�,��Jfi!P� ��'' mI��۵� �� P�� �"�"��i�Թ 323F]3��3 �D r	AN2�8D�D#A �qޛG                             L�@���!f�6��Cb�H�"o��)�mi�"�PI"np�!k)p��k��#�i��O��W�"�/�G�&!.J�/��J�
����M"b!Q⠕�Q �o
���I"b!M⠕�L �oK���G ���F �oI��� G�bG! /���!!B! �������   � � �	7
�J� ��	�
t��� �,�Tb
�o��&	6� �i\�]��g���$樝{� @��˸&� ����BH��ͩ�   ���H�� ĩ���K��b(�ͨ� �� ���D��b@
�
�Q&�/R"�k ��&!��,�,�+!�l!t=��!�z�<"�i;)�f��H/ �F bG� bDQ&��bLQ bJ� � � /�i�e:�(��g����Kie�C(/�g���������$� ����I�� �ʠ�̭ˠ��K� �+� ���*� ���� ��*��+�� ����ӽ�� �������(����A�o �4i)3�&���2�r�� 71� �fj]�b`�\g���� �M&jiie�: /�b�`d�g��h��� ��O�fji�e:� ��b`�dg��h���� �Rbjibe�`\�g��e��67f_g���� �M&R&ji�eb��:� ��`^�_d�gΚh͚� ��O�Rbjiib�e��: /�`�^_�dg��h��ݫ��&�@���E��� 0�H> �M&R&ji�be��:� ��`d�g��e��C(/^d�g��e��C(/_d�g��h��� ��O�Rbjiib�e��: /�`�dg��e��C�(^�dg��e��C�(_�dg��h���� ���'��'����Ձl�&��m��� �� �qr�^T�`�	B0LT"``n�Rqq���
��(��H��^� ��/�M�O�Rbjibi�e6�<7b=dig���$�ie��:⠩�<%&=&&`��%<&&=&dg����$(/�e�:(/�g��i�eC�(^�dg��i�eC����8!.6�/�9�!7���8%&9&&�/�6�87b98d9�_��%8&&9&dg��e��8�!6� ��9!.7�/�g��h�����R�����@L@@F��D j	R&O&���`��$ /a��6�&7�&6b!F� b��$�ie�C /�6��8&7�"9dig��ie�C /�8�%9b&b���68&79&8O9_I�%�8&b9dig��h��i�e��6!.8�/�7�!9�$�gȚ�$� ��h��� �   d��� i	eߒ(��m��m	������(��m �m	�����g��䫵�DPx鄣��&��\i���H�f��]i#ob`��/�^�_̝G���� ����6�/�7����#�/����)R bQI �Y�(Z�!�bK���D���bbY�/��!�;&F.�&6<&7=&�_���Ur�k��R  �ߴ��
{�/�{��&,���   ���7-� ��-�խ��݅խ�-;�-X�-�&��-V"����Ι(��vY�����G�/��5���&.UBb ��G"�a��O����G"�a����[N� (�E("���S'&'�J(�J�˺�/��G�/b˛s�G"�-�����m��lp�;!.k��R��� ��U&�GР�����@�� "b���"7�    ��&��Ȧ�����-�խ��ݏխ�-;�-X�-�&��-�Ο(�!viu*�ȩ�U&�t����m��l�m"�*G ����-ž��w�u��@@�L�� 67���(��;;&;@/�Z�����Y�����O(�ܻlR;$f�*�6���ת�x�f&x�8xkBfxc�i�i�J� �U�� �� ����                                                                                                                                                                                                �,   ��@�.��                                 ��"   LG�2                                  ��"� P�D ���2 @����ͻ                                                                         �6�/�7����>&W)&Ҍڀ����Ԓڀ���->�-X�-�&��-�Σ(��v�u*�H��G��� ��c��6!.8 /�7�!9� ���I� ��c��6!.8 /�7�!9� ��� �[N� (�(E"���S'&'�J(�J�@�t�O���*J.���m@��m�0l�p>�!k����                 	D)"���*J.��K��@�?�B�Nc��M(���W)&*G  ��6!.8�/�7�!9�(������)��A����̨��X� �>�&6O7B(��>>&>@/�Z�����Y����>�k ��խ����-��-w̛ � �>�n66&6.���7 /�6���7�k@��� � O�E�*� �!���� .!6O7mI��Ƞ:�l� �
.
��m �-k)V&-�	&

d	6(/�q�m�
o)p�k
��J5(/�m�5�k��cm�Omّ�Ȼ�� H��mX�Bk)m��Ak)m��@k)m��?k)�C� �5�������i,��s��(�� ��j�(�� ���� D����� ���+ 	 ��F�J���s� � J'b�op�o)p�
�o�D��'���(6�)7

�D������"�  � `�mi ������̞�̬�������� �,�Tb	g	�J� ����pΝ�p����pɝ�p����p6��7��	�� ��6�87b9<b6=b76b���7�/�\��ҽ�խ8!.6�-�-�����-wכ@�� �`b�� ���6��6��&��&��C��F��4�@n��"�n��"����F��&�����"n����J������             �����Ϝ��������5��ʸ��Ш������U�ҭ�խ��-�-�����-w���@��խ�����-wڛ �/@ ���ڀ��������������-������@�(Rxp@  ���"��&���S�*�0��!<�-]���4��"D���*��C���*�  ��

b	t�����*������*(���&�h	t���[��(��	t���[��	tĀ�����(�b��� �� �� �� �� � @    �
���
�b
c	t���J蔫��n������� ��@     ���> �| � �  ��	&X&� �����
&�&W&
�6�'	O�������q ����� �� �� �� ������Ԡ/�֢��bD�����#��r����F�+�c��c���aG����>!$ �
 ������ ����*�&,!��"���?����� �k�]O"�62 ���6 ����� ���b�Ȃ

�
���
.��ț(� �F�n�� �Pn)Pn)Pn)� ���f��&ô&��@���/�O�����"n��ɴdʳJ�Ĳ�����    ? �� �� ��� ��&�6�
.

�����֊   �(в@���/Pn)� �&��!��"�� ��n)�n)��	�8 q	rҕT`!�T@SX��C ��ـ �qr�N �8P@	���� r	 2�0 �� �r �5v� � r	 8�0 �� �r�� D � r	Ԅ  @� �r��`3 � r	 2� IӀ�; r	 4�0 �A 6� �r �21��IӠ5X� � r	 2�1��A 6XN  慰��HG1L*�����D q	rҕT`!R��@O� �r��υ� AT � �qr��DNN �P �� r	R���T%� =	ES��K q	r��DU�RA��D����� q	r��DT` R��O���� �qr��D@S���K q	r��D��C� @� ���TO�#� DT � � 0�� �   �P����� D q	r����4υ��@} � �qr�����4 � q	r�X��4TS@�� q	rϐD8N�P��4TS��� ՁC�N� q)� �qr��C���E� @� �qr��C�S q	r� T T�A��4��E��4��; r	��2 � q	r�� H� �qr��TR`P 0��� q	r��DM T� �qr�� E�D�O1C��1N�� q��@`����  ���ߨX�è��S�  P�ӈLC Q�T�A��8�S�� @   � �ぁ SR�� @� �  �   � p� p�ԃ ��!�Ԉ�z� ��L@8� ���X�N`!TԀ;����TX�	3� ;                                                                                                                                                                                                