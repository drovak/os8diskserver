����  � �  ?   -   ?   ?  	 -   0 ���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��������?�����������(��� ��(���c��ǒ � ��έ����D��DơJ��,ح� ���į����������<��(��(��̀�� ��ά���� �                                                                   0PN6Q ��
� ���,�����������,��������������,��������́����,��������́����,�����,��,��,��쀀�Ԇ����!����aƮ�ӵ�Ӿ��Ł�!����ȡ�a��!�E��M��C�D+�E��F�Gk�����k�+����ػ��+� �             c D��@  ��� ����׀������
����
����������������������������������s��C��EƼF��s��ɼ�μ � �����������������������������C��E�������� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ^^��R1 S� SRQS���AR�a^                     ��w��w��#��7�^�אq�~��w�/��Nr�x��w�/@�q�/~ �7�r�ǐq�/~@��/@�0ܞ�w��}���^Ö�`uT	�� 6� �ՓgN�!��wMN5CT O�#��5@xՓgN�!��wN%��G��t��w^����rL� �����; ����� ނRI-r\ ��p��  ���wMA���^yPV`�L<Ҟ҃L�%�Gyp΀���w�^}����~����~Ӟ��	s�x;��ɞ��~̞��r|��w�~Ş��~�����}��w��|�w��r׀3�q�^}��w���q�/~��GN� x���q�/~@�'�/ �q�r|��w�/@�q�/~@�w[��Cq�Tp@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ^��L`!��w�%5��^�#LD̓A�3�hy��w�C1	�S���$ � H��w��4-�7ހ���E�H��7e��       �^��	8�1��PM�@�S��!@8�^��C�ɇCL�@�^��	8��18M@��w�VN�!���瓅w�N2���>���L`�E8Ne Ra��D^ޔPT�DA̓A�3�R@ze��s��0�z��4O5S�iS%��N ��M�%h�CqI�V��(��E3���N��8�5��D1e��TV�L�#nX1��wNS"((ŖDRe�	v(XX�D	�SS�iS%��L(�S(S��e^^��P@`�RC �T ^��Y!�R  N ER��@I�^���0`L� 2�H %��DO�#S(NS" !�^���0`ÃT`���w��tT^+                            ��CAI�I��4��^��	8��4�VDL`!�E3��w�Bp8��4�V``�#�4��Ҁ7�^���0`C�I�-	��F5��N 	���`�dC@^��M�`	�	8�T5���e8��^�S�`XCI�XTS T�T��^�S�`XN `	���@�`6R���O^�S�`XN `��3�RA��D�^���0`N� �^�S�`XCI�-XT�`R��D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �       ~     - #  1                                �+�� �        �� 	�3!I�!       ���o ``� 
 9���"IH�3 �9�3��@  ������`�R� ? ����Ef �~�	~�/���&��)���i���(����~ ��~�	�� ���6��C��t��&��'�b}|��sH����&��7��TұJ�����3�{9��t%z"(����t���& N� �    ������(�������������kȀ�� ����΀�� ��0NW  ���#����� \ �M M	��À�O�K���4(����h � ��b?yb@�k ��?&�@&� ��4b��g��D���    ���4��c!x� ��� �	�̦&�'��B��t���!�"!�����ζ���K   ���k ��
.

���}|� �                                        �\5+�Ad� ��w���/���� ������b��7�v"�����$� � �v�&����w�b��K�u� t���� �䜴����  ���E�+ �v�&�B�������	����r��޺괾餾��� ����������H�����,�n �������� �                     8( � B6���O                                                                                                                                           � �/���z������/���!&���&�*��+�q"w�� �          � p	��o) ���d� ��o��CH��z�/������ ��o��CH��z�/������ ���cȮ���J��+   ��b�Ҋ�&�&�!>ߠ?�ޢ!�����D�ߢ����c�d��N�+��B�߲����ߨ?Ӹ�      �4b��c��t�2D��                            � ��p)�����f�.&/�b��c(����/����NI��J��2�����B�����&���9�b��K��� �   ���f��f (��&��6��C��ly
�    ���$� � ���&׊,y� ��N�+&� � n	�&Jm�GI	f�J��+��KYfNb F � �             
	�.�?�0� �54&�Q)�p)���5.&/�b�6f���H���(/���������5�"./f�泱�H��z�/����������+      ��9���(/������6}BN������6�}N)��D����њ������� ���6��C��dJ � I	�����K�J�Y��Y0� 0                  ��`���� ���i�(/��������"����"@z���'��N�rm�����~	������/�����&��rm|�m��m���l�m��   }��/�/o�Ƣ�.�.��.'.�K    ���0&1�b��f��&�����c��

�
��}@�Oi�(/�}�!������J��K             ���)`��	���� �� ��i���k�&�����s�!.��d�����t������{)!�������/�����J�j+�/��������� �      ~��A�i~�	��� �L6�~	�� �                                                                                 V�X�ߟ�� n	�&-&-h)�-��5&-g)�-�-p)��-9bf���3f�����'��)�����F���6�/�Ƣ����-��d� ����x5����9�W�u��ߚ�ښ�Ԛ" �          �3Ji�B�I� � �} |�&��"�{)�%bz(/���Mi���#  N   �                 ptHP n	�&-&-h)�p�����o)��-�n-v�J) R I��T�������-B�k�e�d������+E�S�N�   n��b--bhʚp��-�K����Z�͚�-B�k��Ⳁ��S��BP�BP� P                                                         *9 ` �	:�ly�Ji�Y�I��d��J��YI	~�:�����ᘐ:����k�2H����&����5&�g)���9<&<f)����<b�y�   ��7&�.8:d�c�5�b~�bL�p~Y	��:�/�a�ᐊ:�/a �J��YI	 ��d�� �J��BI	 �x��(�� �                  GH�6�Ͽ�hDZNBTFE_ N F`E`_ `�ۙ�E��t��Q��a��L�   �������� ���b�@.�/��N��+   ��b�@.`/��N��+   k�2��g��&�(?�!�&�/�ߢ����ߢ����c9�ٺ�����J��K    �6�D(?�����6�+               �6���� (���+��  P����76�
&
(?�˦
�6
�6
�6�����f��&�
� d��J
(?�ʦ�������8&�b)��J���
�!7�7�e���� σ��� �                                                                                     UGKGU ��7��+i�  ���&��h�������/���8�J� ����_D�.���8�K �X�=u(��^s ��D�򲨱���&� �H��=��� ���N��ˀ7���g��&���&��H��x�_��r

�_���7��B��/́�8O�+�� � �
��T� �                � { =ȍ�u"����^c)�����/�<��y�H ��:F�� 3����(&�%&�&&�!&�i�J�pFPI������~l�Lp�~	�����K �	���к���J� D I�~�ʾ���2���J �DI	��J�]��Z������K                         M�6�N�~# -1  ��YANM Y ]N�Z �Y4N1 Y 4 � J	�S�I���������3�d�Y��N�� � �4�bQk���"`���!.2�bP�����" ��]јZ  ��������]��B �:�a����jD�� �                                                     �L��6�
��!�  ����4Fm�(� � ����44�b��� �4�&��4H��������� �   �1�10c��

�
�0}@� �(|�|} |�'��K   01f��&��&O ��ф������Oi ����J��� �                                                               .�p�Q �m�&��6�>B\�&���

�
���Õʄ� ��}�(����b�(/�l�����| ���ɵ)�[��`��>�����!.��&� �����b� ���bz�/�~�"q��m)� �                                                                               ��� n	~�Ai)~(�~4�~2��Ab��i�C�(D�����������/������������w !���/��xb�����A�/������/�����Śl�)� n���������� ��������͚�!>�?�C����~��D�/�~����CK
cK
 9
      �    ���៫�%�����º غ]Ż �!�⨑���&���wZ��l�<����K �����ǁ���w Z�&�!.��/C�K� ���H�CO�s��Bb����w Y(/�t�����+��槧K ��!.��"�����)�«�,��|���wX��k ��!.�w ���� ���/���!������Á��ၾ�w X�&� �             � �!�⨢���&���w��l�<�Bb����F⠠��!.�\ ����F��/�� �������|���w���b!��(D���\\ �B��F�/F�K ��HD���s�B�/��wY(��t�/���ؾE�d� �WG&WH&��&��&EFfD�k                                 �G!.HE"�����)�����,G�|�G�wWG�k �G!.Hw ���� �FD.����/t�)��FEb���G!.H�/���H�<����H�wWH�k !�&���N� �X�'X�'Z�'Z�'�Cv� �r�	���Ԁ�����K                                        �
�������CO NN EC T� F�IN IS H�XE0XI T�S�EN D� GPET ���RE CE IV E��HPEL P���O                                                                                                                                                                                                                                                                                                  ~/  @ -# N1    � � �(/��� �(����(�|���l���� ��b��� �(���(/��(����/�����/������@���(���j ���w��n�/?��+ ��������(ƚ��\ ��	��(/�b���&� �!��&����K��(y� ���(����� �      ^C �OP �������&�y'����"���݀~�~Ie~I�~I�~I\�BF����&~ �~ ��~�g~I	~� ~I��BF���b�3��F.��"�b�3����y��w��U��"�����"���Y �^ Ν�J_�ʠ�l�Y������ˠ�b��j ��	6܉L	7��J���            y�@�*":=fA������O�"D� � � �&� &� &��⨜���⠾���⨧��w�y��ｿ����a������(���(/�����������/����������                                                                                  ������?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                