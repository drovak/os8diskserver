����  �C �  !< 
8!';
9?>(*%8';% : ';?7> 
 
';?6> : 54?3>(982?1> ;(8';;?';;?> 

0:?';	/? : .;/>(+ 

< 
>(-,+*/).y): )*3?<!>% > ! !??                                                                                                                                                                                                �������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ ����D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �� �  �����}���v	P�n�_��Fn n�&J.
�����ȳ��������R.�i���b!�⨫�Ȁ����}�� %0����&W ��&�@�|"���J"��&���|����/�C��J��B(���}Ɉ � ���k   ? �������������������������������HB�?������� �/ �� R�` VV�!�ڠ/�F����ڶ��r��x|b�i�(��m�������(��m(/�@��|��i�����m(/��������z�� �"�b� �F.��+�(/���H��bV�������m /���ڨ/��� ����� ��c�(�������F�� ���-�����?8��W��2d�pD�F�&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{ �(?��B6� � �gWq���� g�t��D����/���}�� $����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ���������  @��    �bH�
��bmF��B@���Pn�����彀�O��O��������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�׷�����2X��(?�
�

��������������o��R1��D��� N E��D� �@C� ����	��T P�ل�MA	O���� 0���/a� �&�	&�	��J�g�v ��V���T� � � �? ����   � �;: .!/7;?  ({;5(6 (5 | : : : : : : : : : :  	   	   	  	       	   �����6��6���H ��� >Р�����c�c��{0(����bm�/mm"��bm�&��B�f��Ɉ ����k�c�� �������r`���O�֮��&���Γj � �w�?���&��&���?r��/�V��/����yN� PT0B# �텿��f����dw��DW�b��f�Dd#pD0 �TE�RM�IN�AL� T�EST"
DfIKiLAOB.�SV"	-�08/-D�IK�LA.-Bb		�KL�8-$JA� L"OO�P bBA�CK+ T ES T 
D!IK?LB�A.�SV&	-&08&-D&IK?LB/-A.		bKLl8-�JA  T�EL'ET�YP E TE/ST�
/#D�IL/AB�C.�SV!	-.08!-DIL�AB�-C			LA�36�/L	A3�5 �TEfRMbINnALf T�ES�T/
#�DIbLA/CB/.S�V	�-0)8-�DI LAbC-/B	�	L�A1b80� P7RIJNT/ERK DBIAjGN�OSTI/C�
D�IL"PA�C.�SV/	-�08�-D�ILPA"-C�		.LE&8//LP�08t L�IN�E �PR&IN�TE�R "TE�ST?
�DIhLP�EAh.S�V	h-0�8-)DI�LP9E-�A	�	L�P0)5 �LI NEK P�RI+NT ER� T�ES�T
#�DI�RX�AC�.SV	-0�8-DI/RX�A-/C	�	RbX0c1 �FL�OP�PY� D�IA�GN�OS6TI&C9
# DI
RXCBD�.S�V	�-0�8-DI�RX�B-�D	D	R�X0 1 �FL?OP�PY� RDEL�IA�BI?LI?TY�
�DI�TC�AA".S�V	�-0�8-iDI�TC�A-cA	/	T?CO�1 BATSI�C JEX�ER�CISE�Rx
#DJ&CL(AA�.S.V	o-0N8-�DJ�CL.A-A	{	O�PT�IO�N .TE/STK 1� A�ND& 2&
t#D�JE�XC/A.�SV�	-/08�-D�JE�XC�-A�		(4-�32�K <PR�OCES�SO&R �EX�ER�CISE|R"
#�DJkKK!BA).S'V	�-0�8-�DJ�KKB- A	�	P�DP�8/A CPU 6TE�ST�
�EU�ZC.SV	.	-�08�-E�UZ C	�	T D8(E �DE(CT(AP(E /FO�RM�AT�TER �PRoOG)RA"M�
U.DTkFA"A.�SV,	-/08�-U�DT*FA�-A�		&TC�01c/TFU5�5 �DE�C �TAPE� F�OR�MA TT(ER(
�UT�DEA.SV�	- 08-U�TD�EA�		�TD68E) D�EC�TA)PE� C�OPcY bPR�OG)RA)M)
D�0A	B.�SV			�-8	E-�D07AB7		7IN4STTRUDCTDION  TE 8E -D"2C`A	�	P�C8�E �HIg S�PE�ED� REA�DE�R/ PUNC�H �TE.ST/
�2C�A.JSV�		�-8�E-D2&CA
		�PC�8E� H�I xSP�EE�D �RE�AD�ER/P UN�CH/ T�ES�T�
-"D2&CA
		�PC�8E� H�I xSP�EE�D �RE�AD�ER/P UN�CH/ T�ES�T�
O&N/COF�F�
D)2C�A.JSV�		�-8�E-D2&CA
		�PC�8E� H�I xSP�EE�D �RE�AD�ER/P UN�CH/ T�ES�T�

"D2�CAD.S�V	�	-�8E -D"2C`A	�	P�C8�E �HIg S�PE�ED� REA�DE�R/ PUNC�H �TE.ST/
�8E -D"2C`A	�	P�C8�E �HIg S�PE�ED� REA�DE�R/ PUNC�H �TE.ST/
�F�
D)2C�A.JSV�		�-8�E-D2&CA
		�PC�8E� H�I xSP�EE�D �RE�AD�ER/P UN�CH/ T�ES�T�
A*		�PC�8E� H�I xSP�EE�D �RE�AD�ER/P UN�CH/ T�ES�T�
�" ���� � (����B���ǉ�� ��������9���������>���������ɀ 5���K(����� 5����� ���s!� ���)��)��F������< ����?���f�i�/��́���3���&��J�* �	G �偼�|�Y��`��ˌF��:�?߇( �UN�<1��?  �i	 �;`.  � ���/        ��                               0S�E�����Gf,v�Ε��U��U��U��U��U��UV5 y)H�P��� �`��wD� 
   ! -/ 0: ?@ \ �� �  �/��������������������������D򈋪��(?�~������&���lZ��EQ�h!Vb�/�g��/���*f()fU&eF)9A��>����++b���1����-Ι��&�/�+��6�7����Qi��7�8"!!ch��""k ��/��҄�� ������&��J��J� ��3�
  �bD�.Hs�b �J��"�*n &� �|�-��/4��e�FN�B��3��-��/�4��eF)NB��3��
-/4��e�FN�B���'��e�FN��3��
-К/4�1 �NB��3��
-ݚ/4��e�FN�B��3��
4C�BϚ3��4��e�DN�B��3��
4��eF)���3��N�B��3�	�
4���&;?�C��E�  ���3
�ꀡ�x�`b64���&;?�C��E�  ���E���E�3��4����ebF���B��N;�?��E�  ���E3��
�E�4���&eF)���B��N�;?��E�  ��E�U&5��E3��
2��!ub^b01�-��!��-i -	
/�41�"1��!��1i 1	�!�!!C���1 �5 �P(/i �Oy��m�L'+�b��2 �,�/��ȍ�1i�-i�5-�7-�E-�VQ�f�����&P&,&;?��E�Y́\�bbb.���|B�/�\��j1 � ,B���Qf����|B�/���Z�U&�e�.-�y1�y,����-��1�� O)1�-�1��-��!.O1�-�1��-��5�B6)b6���A&(?�6����2r�bn����.����.)�J1 ��J52�&`.)O�\�.��1�����b\b0��.1�l���&���!���1 �5 �2l�be�/��|�_b.X�.d�.���^.)�J1 ��J52�\&w&0)1 �|B�/�5� ���������=�(�(�P� !��&��X�U* ��OV&H���.�Ow��N��w�����k�ZB�M��Y� �C�A9mHC���|�+��풁��[3��$�#dͥ{n��&�wU���`V�Nt;5�z�x������]�P��7-���J��
)R#A�g	3����R��p�mq�{����Ϥ����p�2�f0�����,��PΠ���K����                                                                                                                                                                                                �<���_�w�j@L��|��sa
�5���8�4��PYC�)q���P	WE��KH��q� 4i��C�F�>]{�������t�k��`�4H��7�� ��[�t��>/��lM���局�)GC�'ř�o�����ԣr���7^]���K�&v�-�q�N!�]搌w�Z�(72��                                                                                                                                                                                                ̘B��O�u>���f�M2ܾld��%pfjPw�D�fIQ;����_�԰*K�F}*G��^H��{�m�;*�%�e"��c#��Z�o΄lyg�x>ǵ8�� 9e�cɥ���A���0����Q'�lk��?� ЋXK�V� Ĺ�V�v>t�$���bҰi!�ڮ{��(�C������OnQ�q+N�                                                                                                                                                                                                 ��M?�`�`<a�^�'������x3�0aJu��
���*�O���>qx�r��˖����K��+-�lPqm�sW��#��W����3���E����W��%�a����oh���t�	N��"��m��ѽ�p��3X���k����f
�)W
IK��.�\���׍?j�?������y^z�Г	A���                                                                                                                                                                                                ���6��uja:��R���Jc���9}���0�V��5I.������ÐE)��\��\��]��Q���U�aQ-��?D���}��O��z�pt�Rt�qu^��6||�=8���S�����BmG�����m}�{G��D�I�+sa�yw"7h�ynt{�Ҹg]�����}A��;�{�>�"T                                                                                                                                                                                                ������!���8R���r��mH��s M�üq(�Sm�J2� 41$}> ��P6�������W�a���h��6xS"����?�@�cw�~�����ym[*G�����S��~n�;B#SiF�茢�Ui��`M
��֖$a8!5���[w��	܏��&i��K"�R��2���ɾ{                                                                                                                                                                                                 ��nbTb!:i�=�e!x!#���t!#���|!#���q!#���è/�d�MÖ!A9>��!D�-�#��-%����&�"ȃ��!�!�b���dM)!M9��� �       �X�J�W� �"�J��"�J�� Ё���U��U��U� P��U��U� P���P#� ��V1x̳�@�����D���� �                     ��"��" �3 ,D��D� �                              � E(?U                  >I�Wf�q���������ۻ����I��C1p-�	� x< �N%�	AG��CB� ����M5�=8 ӊLC U�#H  ��ҥ= � �W= ��TN"�P`a�C@`΃	�Sk ���HM�P� H πN3� @�S� �X  ��  ���#8   Ŏ�8�� H��N %�EA A�L0M�N�!  �TT� 4� E��HMN"�  E�TB�4׃�T0����`IÕ5���T� !�8MN"�VI�k �
��C�D	� @P� 8 	���4I�3,XT�    ȀR�	�3�ή��0��3`�NBL��R = ��T׃R�&T���N�k � ;�T׃R� 0� ;� ENB�TX�	3��:� ;`VD��C �TT� �ˣ ����C`N%�E��	�3�m�m`� 	� 2��E� mmz� � �Q�HE �TB�� 8 N��S&�P��H�8STɅ+R   �����@������3� �@4� n�@6� 7� 8� .�@q� r� t�  ��D@`�d,X�R1�� �D`�,E���R1��N�@�D`�A�H��CR�	3� 0�D@`�d,XPRT� �D`� 5� EF�RA��D�A� ACD�ԃ�RA �D`	 � 5� EF��@R� 1CD�ԃ�RA �D`	 � 5� EF��@R� 1NXQ�@D	�R1�D N�T`��D`�A�H��0D&	΃ �	��R-A�T NB 1�O��N2�T`��D`�,E���DT�	ƃ N%��C �TD@�n�>-)n�J�l�s.i ���z�ks&. ����x�+��k�@o&@))$*�on6oH.���ssbo}rF()>-)�n�oorz.i ���o�j�/�o�����ʋ��_T@ �l!�P@��� D            ��/   	���"�K � �$��2�1L�� @            �k�cn&�+�no&$}�F())�� �ns>b-.� ���o����+��co&� �s$i)V�}()>-). ����o�JGp&� �)>�-.� ���p��n���������kcbn�n+n�o$i?}"F())�� �ns>b-.� ���o��*�ao&� �s)i>-). ����o�JGp&� �)>�-.� ���p��n���Ø���Na��C �D�U �#	�S ��A3�8�8��1�ϋ���8�NB�C�L �Ʌ R� 5L� Q�$ �D��U �#� 0�D�C��3�O��8DVC@��5DC�TɅR��C��R�� 8�(�� ��TO�#) DT � � 0�� �   �P����� D �  ���,��/�ʃ���ړ�-�X����ۣ�������&VV��挌���n��0��&��>�!��d��6��CF�昀B����� ���Ԃ���(��Ó���8@��J��/Ԙ��������b��(�Pn�/��B@���Ⓚ��(��������JX�����/�-��}� �?��}�