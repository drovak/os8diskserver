����  �� @##3	2/  u2> 6 1 *+< ?1? 11 ?2v (���������                                                                                                                                                                                                                                                                                                                           ���6��C��d��6��L��&�� �����   ��l�
�    ���&�����c��c��c��c�(��&��0��'��<���  ���Él��<���   �
��'��'��'��'��'��'� � �         ��D����� � �B��N������I��La݈c�mX��������������� ����l��&��<(������ ���L��<ҡd��N��b�� `� � ����ǉl��������&�F>�����J��C��
��D�����J
�����4�  � �    ���Ɉ� ������ J
�
I���&��&��&�	�t���z�����?[���#�߀���� ] Ϊ^������ ����l��(����� �����"��h�!>�&��<��X �� �� ��������l��˫*�ƺ������7��B

�����'��B��d�� �D���oɩt� �       ��� (��J
�
I��@n��#����툘� ��̲��&��&��&� ���� �o���D�ǫ ��\�W�C?���                                                                                                                                                                                                � �i �8"`7�+    ���/               ��/      � ��r	  @��b("�jb5a�� � �� �?�Ň!��� ���@��� �4!�"�� #��W���`� �/K�"�
�F���� ����V����2�  �����"�/�%[�)!��� � 5�����n�&�&�n@/�������nb�� ������(���H/���@���'D�������(/����n�r�b�b����(��b���bcb���/��"H����)���������n �bD�.@� G P���`�������=�� ���(��(�K�J���������&��(��(�J����"�����(��ɹ�����(���(/����(/���(����(��ɪ������������ �               �&D..��+ ��Л�/sKdB����b���-榣�,p������cH/�F���� ���������� ����� ��                  `` `` `` ``    `` ���             3���33���3��c`�`���g0cc������  @� 		H`` ���1���1`` `` `              0` �� �� �� �� `0 �` 00 00 00 00 `�  cc����?����c<c � ` `` `��`�`` `              ``  @        �� p                     ``   0` ��  6  ���7�3c�Ã����{`� �``` `` `` ��w��� ` � ������  ���8x ؘ�7��  ���  � ���� ����� � ������������0` `` `` `` ����c�6��������������         ``    ``       ``    ``  @    0 �  �00        �� p �� p       �00 0 �    ��0` ``    `` ��7>f~fff~f< f��s`� �l�������������������7 �  �  � ���s�������������  � ��� �  �������  � ��� �  �  ���7�  �����s�����������`` `` `` `` ���    ���s��0���0���  �  �  �  �  ��������c��������c�3�������������������� �  �  �����������������0����� � ���0������`` `` `` `` `` �������������1�` ���c�̛���c���6���1�` `` `` `` ��� 0 �   ������ �� �� �� �� ��   � �1�` 0   �� 00 00 00 00 �� `� �lf```` `` ``   0�  �?� ��0                                                                                                                                                                                                   