����   H t �                                                                                                                                   >                                                                                                                                                                                                                                                                                                                                                                                                                                   �����۟h���!�⨖���b�(/��"��c��ˁ�Ù�����۠n� ���Ȁ�۠/�Ȩ� /��/����b�(/��"!��(��!����bݠz�!,�&������&ȟ� �� ������H?�����ʀ��ރl� �   �f������/�����Ã��         4���� �lܕ��~�3��������#6�"6��Z�?'H/�'����`(滋��/���!���&��&�t�ޤ����l��{��?(�l�!>��?�������#b#b!��"� �b�b%�b&f�bf�'�(���@/���'�b'"@��!'��k                      �� ��R�� {��p�&� %$ !f�b%bb����� .&�"���$&!�/�!��%&�)&�&�')�J&�&�!��� &�!�!.�/����k   �����r��r�{� �                                                                   X�WV�|� 0� �W� %(�/!�/� �!�  bF �FF��+f,�j+!.���+�(�,�+�"+,b��/��� ��&����"@�����	&�)&	!>�?�)��+����,!.)�k��K                                                                            ��w�� ��P�� #f����)����+b!�	�b��I  
  �&�i��))�J�&+"	�f�,"�	�,!.���� ���c��F�)&�)�J��"	b�	&��J� �    ���٢�n�&����Ù���@.�/��J� �                                 �� � � ���r`/6��%�%&�&&f" .&&�&(�/������r&���b�b�i&&���#�&�����Ù����/������(���� �F k G D                                                                             &{�68S���SO � ���D ��Ù����/�����0��ϗ��"����%)���&&�i�%)�%)�"�!⠮��"���%)�&)��;F h G  F a G  J                                                                             �� 0��C�O l�OZ������"������L��(���H/���%��/�����&&&�"ș��&���(��@��(����!T���i޵J��%��(����&�%)ߔ*�*�%)� ����"�����!����&&�j                     ��$[ �?�^� O�� 0_����� ��i���&)�F�"d��/����/��&�%)!.��/���b&�"Ȁ�� � ��&!.H/���n"�b!���g����/�դ�֢�d����b��s�������Ú      !� ��D�!�7������K                       �_6�S �P�  $$s$�@���!�b%�k ��K ���B%�k �b!⠥���&!.�/��������)�"��b�kY     �@����ƶ���c�(O�Ƹ� � !�&��������i���� �                                                      ��  62P�_ ���s(���HN(�������������w��'��������֙<։|��D���c(��*c)c�*ǉ*�)�J��������7��'��������'��'��'��'��'��'�,��r��r��z��'��� �
��ǀ �            �a��ܾ�̦������/l ����`֡��P����E�   ��(��(���������������� ��)���������)���������������'��'��,�|� �&!̯��� �                                                                                              �+p"0�   ���Z                                                                                                                                                                                                  ������W���-��������_��˄  �ev�eW�� �"� �� ���3+24Q9Q�9RK0m����N�oB 
 wx$ B��Vā�������3ԀB�n�$��@�nN� � v �(ǁ(Ā ���l��<v����
�j)                                          ��?�����b��j��b��c�(O�H������������,��r��{  ! �&��Ǿ�'��'������ p�����s�J

����{�P5� �                                                                        l��ր�����@�� �)��C�G��@: ER /S YS :T EC O. IN I/ "S YH XW HK '@ ^U Z� ���MW +0 ES ., .X WM Z^ [0 ,0 XZ ES "N 0E SM X'   @ I� ���@: ER /S YS :T EC O. TE C/ "F ^A Ca n' t  fi nd  S YS :T EC O. TE C 
  'A ., ZX V. ,Z KM V. ,. XV                                                                                                                                                                             *<�Qk�����͙��+�FY�fr�}���Ԫ���*I�`��*����-�?|̞����<�Il le ga l  Co mm an d  @  Un te rm in at ed  C om ma nd  I ll eg al  Q -r eg is te r  Na me  @  I nt er na l  Pu sh  D ow n  Ov er fl ow  S to ra ge  C ap ac it y  Ex ce ed ed  S ea rc h  St ri ng  t oo  L on g  +  Im pr op er  A rg um en ts  I ll eg al  C ha ra ct er  @  i n  Fi le na me  @  n ot  i n  an  I te ra ti on  A tt em pt  t o  Mo ve  P oi nt er  O ff  P ag e  wi th  @  Q -r eg is te r  Me mo ry  O ve rf lo w  Un te rm in at ed  M ac ro  O ut pu t  Er ro r  In pu t  Er ro r  Fi le  E rr or  O ut pu t  Co mm an d  wo ul d  ha ve  O ve rf lo we d  Nu me ri c  Ar gu me nt  t o  Y  Il le ga l  Ch ar ac te r  @  af te r  E  Il le ga l  Ch ar ac te r  @  af te r  "  No  A rg um en t  be fo re  =  N o  Ar gu me nt  b ef or e  @  Se ar ch  f ai le d  +  Ne ga ti ve  o r  Ze ro  A rg um en t  to  @  N eg at iv e  ar gu me nt  t o  ,  Ca se  S up po rt  n ot  I mp le me nt ed 
 	 [ us e  W  fo r  Wa tc h  Co mm an d]  U nd ef in ed  I /O  S wi tc h  Ca nn ot  W ri te  O ut  E rr or  M es sa ge  O ve rl ay  I ll eg al  C ha ra ct er  @  a ft er  F  @  C om ma nd  A bo rt ed  C CL .S V  no t  fo un d  or  E G  ar gu me nt  t oo  b ig  E xe cu ti on  a bo rt ed  C as e  Su pp or t  no t  Im pl em en te d 
	  [u se  E O  fo r  Ve rs io n  nu mb er ]  Un im pl em en te d  ch ar ac te r  @  af te r  E  De le te  t oo  b ig  R ef er en ce  t o  Po in te r  po si ti on  O ff  P ag e  Ex te nd ed  C TR L/ E  ma tc h  co nt ro l  no t  im pl em en te d  No  A rg um en t  Be fo re  ^ _  Un im pl em en te d  Pu sh  o r  Po p  Co mm an d  @  No  F il e  fo r  Ou tp ut  � � � �  � �T N@@Sa��耝                                          ���0J
��❚b��b��h��<��t��D������   ��  @   ��� ���&�����c(���(/���(����)��H� ���)��ß����)������ЁlП8�(O��������� ���8����������_�B�V�� �                � ���i	  �F" =+���� ���&�(?�����O��������bH���@.��/�����������   ��(��(��"�ʊ���D.��&��(��8������� � 


� ���ɽ ��(����������(� ������6��6��C��i��&�(����(�(��� �    � �� ��'��K����>  ?�O@�^< ������   �(���i��)��)��&�J.

��b���h��/�����c(����h!�⠗���J   ���(����)�����M�=
��8���� �����(/�ˢ(��ȼ+ ���þ������J
����0�J.
����D��D��J���   �
�"�bJ
�
!���f�.��j ��   �?/     � �      L	                                  ` �          	  
L	� `                      Q	    GAP8W�XSn5׀T�V�+���t? U s5/V��G�Y�x��w\�Ql_� /  ��������� ?o/ޙ*@ _ ��[�S��"&"!.��/L��Z{�A`i@I�&fIV������b�|b��Q�PM�IޟMn�,�&ᤊ`+��h0�*�S�L�r^c�b��&��&�@?�Ii V	��Ȼ�f� �h���hi��fh��L�z!.�/N��к)(&\){>`�Q{�0�/�@�)�"���*j)�:� � 8�I_�l%� F��(D.��l��(��BF�(�K D��l�m0��F�m0J
�
.
�� �m��v0��'� �����w� ��L!�����Hi��b�H�cx�� ��"�""c� �""t"�"�L�ǁ� ���GГ� �@@�p�����Hi��c��cG����D᫢Gכ DV��(����/�!��D�&��� ������ii�_�1�_$�WL�$Jk_��8��!B�$!.%�/���$�J�B&�$�$o���� �H.�+O1_���aB�BI)�B�(�JP�%'&'�"�L�%&&'%&�&�!$��� &�& n''&&v0�'cm�'�z�B�$&B(/J@�$W)L&�$'&�%�!&���&v0�'cm�'&t'�J'%&�J� � Γ`L�B� �_8�L!��Xi�&��&]��Mv�j���JLc�x�
���!���$�&��ch��!��$v0����$���&% .$�/�$��k�o��J ��$Áv�d����B�b$�jO������ꠀ���JY�����!.$4&�$&I���bIX�Oy��Kyk����!%����/���z��      ��8r"@n�Jޏ&�F.�D.�&�/1��n�.����&ˏ&����K��"�i)��K̒Տ"f�$�� �r@.q�/��K���,�"u�"�b�b��fJk՗
 ��ߗ* !��bH����J� ���ba ��O�@��   �J����Jz%�.Jk -j�j�MP"LN S_ cM���/L � ��   �j)�j)�j)�����{�s�@��oM)*I��耀�������*���"��iA�����q��b��/N��{`9�q��Si 3��3f)(&�3�3:b (�H��:T)֨/͠�(�*�|�QI���R3 n �� ���� ����FH?�q��/����6�H?���������K 11333������8�d�b��D&D�/O���/�_�8L�!��I��D�/���.�RI��D�J�   ;a. �/� �:T)�.�R��C�*IP���&� ���b!a�V�L�����w� ξJJZ��`���&3�* ��$&Ii�$b$f@�WL�`� ����b�b�j�/Lh��!gC�&&X�]y� �
\�R���Ji$�''b�W�����'�<v@�����L�R!.L�/%�/L%�$�ba%�/�=��@�
@"@�z
�
��7i � ����
"��n�&�=&�� ���殲�n&m0cmJ
�J
�� w� ��(���(/���(��.�,3%cm3%3r�%�q�/��*o��J�L�  �8�e���� M	*Gb�s@����j)�}Bj)� ���jnu"�0b����u�`oj)��K��}�� �o ����j)�B~�
j)� �H��3[i�<�('&�<�a3���(��)(&(�"�L�)&&()&(&B!'��� &�&�n((&&T)\њ'(&)!.'�/�'�T\�'�J()&�<�3<'#^)[��0 �X �!]i���n^ (9!.�(f�<&��<((<d<�D���   �;�a ☥� :"TF�F  Q�F $��(��".�L�H �H�H�H^�� �##b[(�:�n<;� � ��c9�9d)L9�tH/*0"9[i����JQ)JP�Q�@H�P�� ���F��6�(?������ `�����-&J �OM�k��KL���Q)��	9��hɂ�f���ck�L����c��bv���b�*���&h � ���J�,b�Y�4!b:(& a.!3&34" ��!�Iݑ�(�Tז�(�3�J� ��$�m�$�|$�KZ��<� 3�O���<�I��� ���V�H��wM	㉛w� w ׁnI���� t@~�}�+(T)Q(�3�JJh��Lg W��iI��I��SI���;Z@��Z�_<�<<7�<�n��7�>�<�� �+Q)0Q)��1��L�O1�f��J ��Ji���I鍰* {����{�`)�T�� $v�M.���?B�J$ N�J�I*�%�+��� fykZ��K#�  "!�9^)J�Q��q�/��{`9�����D$����D 18�o�@��  ! "# $  јo�X���&��&f�n��f]ŚM��9d	L�u�/��H.�bbx���F�����t���/�¦b��(���/X��&�.�:/ ���i��6��N��&�p�  ׊lp�    �
��&�"���׊,p �   �آ��� ����LR&I��L�IN��/�񫯷fUp>:��I�7�s�'&�'Á�����(/���'�b�l�p9  � '&��@8���6��56��s�r�r�r�r��rR�b��s�<���'��'�����7�n=�n�c��s@IiN<t�y�O��J��]��b��/L֒��r��{             ��X�4]D*O��v��w���ߙ��v��vu�����5�,p�� �L�R�lp	�y �k��lI���� �F�bm???t� �43f�!>@4���43d���3�$� ��JO��k �f� ��&� � p��J�����>d��݅�6 �� ��Ѣ
�&��&�?&�>&ǀ�LR&L���K   � � �!��m!X���D.F���P��0��!��!��� �      ��c�$bbqI��$&$&A.I��$!.'&$&$!.&&'&�&��&ŉ��<w�(,��`/�(����(��Pn�(������&瀂�����J��"��ba,� 4�>4������� .*��F.��,�" ���E�D��ba���0�������ns"�k,�) ��� >D@ � 8��?�ѹ����vV� 8 �!p@�((@@  �^��A@Si�R��?Qz��F�8#(�V��R��� @� � �(��""P-�?�?���^����e�?$�^��?�/�!�b>�?�(� ?�o?�o�?$����?f�Q�� ?��~��3�<�ci� � F` � >D�1                                                �J&'eIJ��g�`��U f�  ���I��%d�.�RI�VI��� �%�/ Z���|t���? * 
 /Z	LIJ.�n<<<t<'J �b��@������+   �    *  �   ��� [ �� �g�(' 0��!%���!%⇇K O	b��                                                                                                                   } ~n��
n���	n��G�nn�n�nn����n��o�n �r�Se5�sc�Z5�S�er	PWr�`t�		 		 P�[QP�		 	W		 �R+r�S���	�W&��"��"!�b��"��"��"��"��"��"�)발�\�n TS�a����%P�e���Zm)�6�Q�O5J	��4R�k���=l                                                ��B���[�|��B��r��~a�� �������2��s� ց��.�ೢ&��� ���'8� ��Ԡ/�����t�����"���������M�|�����T�|�3�y��Áp�����"��ٺ��
 0H
�� �\��� �����F�Á(��D��ÁD�� �   �� ����_ lI��s�d9�� ���E�/�m�����l��2�������B���`��e�R������������� `��� ��!�
�����{m�(�́���0p�'� �3�cǹd�6��Cɹd�6�O?�|3�J� �                                                         �ol��P����� ��   "# $ �fY� Ui!��b:(&(T)!3�]��3�/�(��3�-�/�g�y � ��fi�ciMۖ%�
O��O��YY�Io����jAD NE CG LT Fc	M,���کJ���H���F���/��"���ڠ/���   !> <" ^@ 	  EF IN OS _Q UX GM %\ O������c�x�
^�?�_�ַf��f�v��f��f��f��f��f��f��f��f��f�Oi��㨠���&N��L��/�KU>�gٚRW BG kl����d�������Lc�M��vH�M�e�@L��ii���J���U'��NKgy��/���ߨy�(L�� ��K� �=�R> <S U�K�����(��!� &Jk VW�f !  # $�&C ���D.��&��?�x�Q˓�˄��8��0��/��E�/��������0�S��p0��� !.��{w�QS�{�?��� j	��� ��
.

��ʂ���    � (o��(/�x�xoj̛ F��+L�?Nx�Q��;fi OiQL��x�Q�Q)��� ����5l���i(���V�u����B���e�ܢ�v4�����D��u��ά���r��/��������ˎ.� �,�� �L #T�PQ�#�CE@3� CR�F�#�@B�@ DM�CT@S� 5N $��� �@0E� Q� �@1�@5�@4� BP@ �@0�@2I�TS@ ��SF� C@`� ���@2E�W� DC@!��0�@2��3    ! "  $I	��kR!.L�/�z�!.%�/�>� w� >��3&�R)3�J5�"��l6�'�8������6�5�p�� ���������6��'**0��l�6� � �
�%��J�LL�RJk@I�I)��;LL�LIi0��.�QJ���� .Jk .��������Á��L� ���X�R�� 0��w>��5I��X����&��&]��p�(� ��OL����|��K�����/��������n�p�1 �
��'��&�p�  I���à  0��I� 7�
���ZY�! . `)! &fi]ʚ\ƚgy�|Q)�Q)�A�H��`��Z`�{�7{�~�����!.��&��6��; L	rEpn)p� p    iiF�$�Z���1>yـ� ! "#  ����&�J�J .�� .��v��"��c��c(J���d��6��C��d��0����7��D�����7�����       ���������oB  ��Cj	Q��S�jQ��VVQ ��|��^ ���  ���Ѓ    @ ��d0
n�2&2�7J �   ��&XhY ���4�b���2�"���!.on�"�枮2b��d��6a) �(����)X��4&��J�"���      LI2�&������O��n�"2�hl�2dS�J �Fo ����J��JI���(� /�I��!.J��$�H�@.0/JI���* $q%�J��$�v��ڶ�ugu�v� ` ������o�00-	                                                                                                                                                                                                