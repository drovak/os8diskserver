����  @ �Q9991:::1;;;&;6<<< <-<9===="=+=3=;>>	>>>>">'>,>1>5>:>=???????  < 8 4 0 - * ' % "                  
 	 	                    /8'65>(*+*%(+.> '4%(+.8 '9+'3< $>$8+'4+
888888 998+'7+$$>6$>*<'2=	**C2  =
8
$
 $?4/?
D </?'><(/?9'=  �+&@ٔ�MA         L �          � �                                  ��    � ���Ѝ��#5�T B�l@./d�f��"U� .P�ZJZ�YZO �dFF�~ .�lBBK�s�
��� �v���? ���?������Y� >  ��&��f�	&f"f�#�$�b�bg�J!ff> �O��>��������������y��/���%�(+".�/�%�(+f.d ��ǚ� �b>$��������� �T�P��Jb&��>6�>)*D���	&�J�u�|) �3�T/��"֕"$����"O���(���bH�� ��b��

�
���)��H����O����i������  &�� >i<�B�"�j�I>J��J����� @/H(�� 6�"c "@/���i�*�H/�����b�bc���DD����r�R���%�OC ��Z�O ����_��2!Bt��Br��/�!�!!��&�&4�O�����t�J�&�&4���D�J��T.����ZCȼ�#���!�B�"T��2@���!⠩���%�)(�)+�).�)% /%&( /(&+ /+&. /.&!.��

�
���&����������? �0�%�T (��@��!��n� ����U�1�2��3&� ��1D�2�������4O2�I�� �
��B1�b��b5�j2�O������5c�J
6�

�5�J5�065d5�0�(/���� ���&�3Á(�͊��� �3�� �Z.
4�33C���32F�1���KD.!�`������ ����f�� ���/��� ���b(����@?���6 �������� ��&�&t��� ��@.�/���"f �d��������� �	��b� /�(/��@�␹�	'	�"����	&�"����+�� �	&	7�'��ؕ����&윿��0�`���@��v�� �/S@8��QCO�3 ����(����bc��!	⨀��J��� ��$�#��#� F��#�|$!.$�k D��b��bb��������    (���&�(�����ʘ������ (?�P�/���J���+�����   �&��4D�$�߫� 	A�� �
��)��/Z�0�?���?��� ���@��o���
��� ���(� ���(��(� �!��&�Ι���&�&�&�������c��b��r��r��{�ϑÁ��J�B�Ȫ�Т��r��r��{�<���ǁ��    � (������0b��)!.�k��d͊��� 08 � �  ��?���������� _
0F��]��_��*��'��,��s��v��E��\��9��<��-��/��=��3��>��M�� �E��s�� � C �X�,��Sl�R� �^)�]%�_$�U-�S.�T9�E6�s6�W2� �T9�E9�s9� �              !# %& (�
��(��"b�'d���?��"�'���t#&#p)|�/!wy�V�p(�                                                                                                                                                                                                f�&�	�Xn�~	�|�b�B���w��B�}H���
���&6B��� D��kBځ�'�~Bxj})���BB�F.��bfb���@�&�&�J� �  b  b �jD.b��B�J"bb#'"+!.!�k��ǎ N� N��J�������@	�('�&6B�F�N}i&7� ��H��ct���BF���B��!.	� �������������
�s�ǁ  ��&� �             �� z� ����5L�p@�� ��5L��@�� ��5L�q@��  �5L��@��  ��� ���)H@� �/�wW?�B��}F��}i&!.AbfBn���@&B:���Bȅ�&&&D.b��J� ��&�� �o� �.b�J `�+�&�� ��$��b�B�����k ��Á����  �������+o ��|��ڶ�g�Cq�T�?(8��_B��!/ a.$/�!�$a.(/�!�(a.,/�!�,a. b(/� �A�$�(/�$�A#�(�(/�(�A'�,�(/�,�A+�A�)b@�o O� �B�-�")H/P@�@���!|�Bh�2�A���k�-&BH�	&)�,7)�,%%&�� �j"$&�&�(�j*,&��� p ���%)"�D.�,	|rA� �	�)�	�|%-f��!	�{� �B�����/���� ���N0�"�>4�E�f1�w'��g���têV��ػĹ����:b݇�����
&�AZ�q��������� -�9D�NX�bk�s{�����������������������������@�<8 40 -* '% "         
 		                  *�U��U��U��U_ VQXfX�eQ�e��UQ�e��UQ�e��U��U��U��U��U��U��U��_��"!F)�/]\���j��Km��e�`��
�
�t�����`g��o 