����    �* . *	 /	  /  /  </* $.   .  $	  $  . *	???.*/  $  $
  $  $ $ $  &���������                                                                                                                                                                                                                                        �h��                � �� � +#�����0      ,~�/%˃}�Z P       �  ���`.�Q�� ���� �� '� � �� �� ���R�q�^ "
����x�"� ���t� yrt/�n�~w�x��n��" �p �rs�o��}�� � ���� �bHN��4�o���F����0�������{ ��b�J H��4��c��

�
����+ �(��H����+ ���� ���� � �#��� �����/��N&Ɂ�	 6 " u���" u��� !.�/� � ��/��  ��/��K ����@ ���?� �s� ���c�(O�Ϧ��0σzi�y�����Ѐc��b�c�(O�϶�>����.��c
�� ��f����Ѥ����c� ��d������Ԣ�j ���I !�i��r����k          	�y����ϳ���ϲ�� ��ϳ����s����{�_�(��^(/�]� �� �� �@ ����8����8���� �b��n&��������r���)��z�)��r�k ��4��y�Ǫ!)���!�� ���4ɴc��F��4�@O�Ȣ���ʴ6���    �
|UY�Ɗ W鎁�|�<|�?SR� �|Q7�|�Qr�jX�U��ڋ�J�S�PO)� ������ |Qc�sP ��i) ���4��n��b��b�b�b�i�y   ��� ���D������B��b��j�J�
��������������)����� ��F��4�b!���"��bi��r(���`/���@���`/���H���������j) �
         胬�Ѱ�/����J��	 &���ª��� ���F��4��b��c��t��D���      �i��h��������&�����������ǉ�����!)�k   ��&�(����(����,�ǚ��h�!)�)�r��/Ѯ������F��!)������������ ���� ������� �� .��d���!)�5�!(��� ������,� ����o����� ���b��l�����<�&6��É�Ϡ����<����ɠ� ���\����<�H�  ��4�b��f� ������!)������hǀ��!)�
�����k 	 �(����B� � ��F��4��h�!���D�ԫ   �n�O�{� �H�/��騻h p � @��
� "$%$ �!��3  ����FJ>

����� ��(���!�� ������纺B��~��r��|��6M� ���F�&����,��|� � ����   �`/��@��� ���b�(/����c��d � �� ���4��b�H/����b�i   ՀN��  �kQ'O#�z��T�	G+�D � ��? �����;�����	�����?��"��ǉ����?���!��#��!���!�������A��������9��!)���!�#�#�2����ǉ���4��"���?���	��#����{�)�>�I��'�\��f������ ڪP�9 	��������������	���!��������!��U���,��|�X���ȳ��!)�>ȱ�#������!������_��!)��'�����Ӛ�)Ӫ��?����r�y����!���'���:X"(������W��`���Q g�3� ������	 	��	�� 	��a��������G����?������#���!)����?��t�f������h��Ⱥ������k�������v����/������&����k��n�p����̚r���{����'� �		a>�/�	�a���	3����1C����ެ��� ���bgׅJ��y������&�� ���"!���!.D���"�i�y����ף��סz��0��'���i� y���i�y����&��0��r�� ��ף����r���0��'ɀ�       ���F ���2�����C�/��<ڻ���������욉 �  �- �KYP�X��������)������>�v������#������p���&��&��"��c�����0(���b!�!���.�i �����!Г����~��!ϒ�!)p�ϠJr��'� �   )����۪�����2������ ����ʀ�`�P� � ��?�:�� �� � R�� �U�����������	���!��������!��U���,��|����ȵ�p��>ȯ�#�������!�����������?���!����!���!����y������2��w�'��� 0��É��c�!ۛ������
!�Ԁ83��:ì@�ڕ�ә 	��	�� 	������������?����������p��>����h���?������#��������?������p�������p����������������'��'���!��S��������y�?���!���o���� �8 ��Ƥ��0��գ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �Ι� �� ��ә�י 
���ޙ �	���� �������� �� ��@���D�0�	3�@�C�U�M�`
�� N$ P�5TP�S         ��         	�4         MG@         	�R @ `                                  @ `      P       �   �   P       � 0 0 �  0 �$� 0                                                                                                          41 �TVU��U2=�C �U��U��U[iiiKCT�Qs� ("(("FR�QT�s ����'*�D`e��f �F))3))3�Ļ���ڻ�Իɖ�LD�O�#/ �ɖ�LDL�`�CFCT O�#` �߃� 	3�8�8��1 � � �P�� pT� �ē��{P��tǂ;|  �����q#8���Tn ����X� �� ��C�l� � : [� ���P�'�|��:�y��7��@�4������p:�Wē�t�� � �������� �� p� �� p �� �ē�t�� p� ��q�[o��� ��t� ��4ǁ4`5N��y� 0�t��� p���1��J���1��JNO �k � � /_�:��V` �N XS�C  ғNP �ԃ�JL�/�� ē 
	� 0ǔ 	C��� N P                                        	� �@ٔ�MA       9 %� �#+�A�                                   � �� � 000D00D00D0:K� C   ����� S�O�^�UB��� R@� � ����dB� ��(�?��s�@: ��M��8m�e��a��$���g2�� ��`���f��?�&O������&��  �&�����1�(��'c(9�(c)c*c+�b��c��|��'��&'�,�8Z�/&'�,�(  7��	�&�l��''� ��s���(��F����" �k�����!�⠺�����u���F.������r��/��朂� bx�/ �"�@�O���U�O�(������'��'��'��'�����r��s��ˢ��r��r�|��'��'��'��'������"�����0�����'��'�*��'��'��'��7��'ف|-�n.�c��r�b�n#f�ɺ�2�dt�q�2c���T��Ԁ8��`e��D�[�̀����/
 ��u&�6����{@d!�x�)�9����
6
	&�&%f
6� D�F.�b(�����`���H/���	%t�J��� ���ɧ ���� �
�<� ���l��&��ó�F��'��+    +�w��n 6��+�(��+d_2(���(/������� ��
&
(?�(�`�z�����b(bi(l�4�lv	�?����2�	 G�� ��7B ��"$� �7�".d�,�����&�
&��ھÈ�ߤ������
��J��ڼ�ڼ�3
��
&�&�
#����J���
�d� �.�n,�kÒ� ���&� �������/��������)�&������(���¨���������b
�j��� � ��t�O\�'e���;�t�����6ؿ�
6
6�&�&!�bc!DN���J�J����������J!�"���-���� �!&(?���"(����/���
c ���J�������"����&�
&�����F.���.pX(ٔ�ȫ    )(�����:X"(������W��`����7W)V��7� 6x���� �3$�?�� �������J>

����� ��(���(��H���)� ��&����k 	7%2 ��	&O�	���%�/��� ��z�.�����fai�0�0/d$�J �       � �� �� �� ֱ �� �� �� JU L� �� �� �� Š  /��xR()\()0�  +t��@@��?���$f�&
(?���(���)�������������$�j�J  �O�����"�/#�K 	��6�� ��/䪤�.��D���.��&�.��(��D��������H.��&�?�
�

��(������(/������"�� �   sn rl sr sj o� � �?0������� ��� ����⪩b�Ī��t�
.
�Ī�t�/�� � 6
��B�b�d��T���� �   ��b��5֢��/����!�$%f���-�J�&���� ��!���&d������&'b��   4
�!.�����7����\�"�"։lց<$���;�/A��!@��������, �0s������&�&#b�b�h�&�&�/����i�����( 2
��&����   	�Cf"H��F��� /������B�� �� �&!���������*���0D.�&60�i6���/�ⲲP��_"���e�*��~,�(/��lr����$t	c%����s���207+�D���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            � �$�Nq � 0R�	�R1��D D�`1����CP�`���sT� E��ɉD��� �Q R��NR��� NQ�T���sTU����7�σG���p� 5��`��7��	���D@RC�R��P`a�C@`΃	�Sn��T�ȓ�X�8��4�-HN���N"�Ss� `���OB��<� p   I�pV�pd�pm�pt�p{�p�hr����p�������U#d�/���"h9�t����F`   �'9�3�� �      ��a�?� ͏"�B� �  0��@�� � I�	E�O2��0N� N ��`1��� 0� �Հ@F  N$ NR E�	�4 � `� 1NB TN %􀎅D@ ���C@���1��A PF(� 0 5	�3T P��5� 0��C� 0�R1@6�DC@N�T� P�AC� @�E� @��E �� 0��`�u @�O3�0�GB�0�4X C �$�  �	�S@�0T�@ T@ L  0FN`� 0��  UVBLN�  �A 5� P	�GR  U�  A WN !B�TEN@!� MN!��C  Ռ0`CSO�#�L�@Ra� 3N�O�	0��C2L  A TR�0 T� PL�P.�VX�^Z�jA�Eu�&�R1�4�6>�bn�rf��xG�	!�I��$x�������������ǈ�Έ�Ո�����������    ����������)���I�  � �
��'�b(lb�v�A�)b���"P�U���k꠹��D��E�S����7RK�"�&�p2                                                                                                                                                                                                