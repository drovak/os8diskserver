����   �������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                         G�i� �;`.:" � ���/    8 � @����  D  h  ����p?� >                           J�7����_nf.@a�Ј �U���? +�G�U�&�� 6��T�o[����f6 @     �x��TGV[ �       �	h��    �� ��J�P��po�r���:o�;�P�!�/�^�������������������bW���������� )"� #��3� 4 E� xV�[,(��x�(w�v(/�u�(��t�/s��r��q�q'�!�s��&sK�*!��"��*p'+o',�+ ���f�h���n �bD�.Hs�b �J��"�*n &��,�m����#�b^����S-6TS'�-1l1�J1�J1�JL��� .11d�m�S1v1ģ��R�-S'Q� &fjb�nfi � h" j�(s�g�/cne bd�m�I���I!��"�����J��e�c� ˠ�s�c�*���/�-��b�p�   �
�@.b/�F�u��#��r���"�a����N���N��N�Q������� N���� �+ NQ��� ��6&�- N�� � NQ������ �N_�C ~B2v ����2�����2��N� N�B ?NC�!z� ��Q���z6&C56N̚ ��7&H֛�R�Tٚ! �s�g"�n�bQF�u�7� �P(/i �Oy��m�L#� ٔC����ؠ�38f44d4!.#�/������D������5�4!.5�/���Q �)/���74b6Hi�����݁�ؠ3�48f44B!(�����߸E���߼������5֠5�55b!4����Q�)�"���7&46&H�� ��������ث��&69����B��N��JB6)b6���A&(?�6���� }	Q�� # �3zg84f4!.#�/�D����z_ 4䌆� �38f4�n4!.#�/�E���ڀ4�!|㠱�4�J���!.tEi��ڀ4�!|���t�J���4�6|c5�h��7Hi�̳�̃�e@���?��b

�
���(� �e(�>�e>�ߋ ���������=�(�(�P� !��&��<���k����q n38fqH.8n4qbzDy���qH.8n(4&D�����q!.�/�q��q�8b 3�qH.8n(4&E�����_&q'qqB{rc5_b		c66b!5���56	666!.5�/� �!.q�/�Q� �3���7&H��ؠ��?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0�H>�%�2�m��ݠ3�?�*8�?�4�h?z'D���E���ڀz�6|c56b!5⠯�2�JQ��� 0?J. �?�@�K���� 3�82f"4&D���(�4�m���D2�Ò��LQ���3�� 3�82f"4&D���(�4�m���E2�ݒ��LQ�� 4��  �������d�� �v �J
�
��(��H����3�8(b42f��݁Dْ�ڠ3�#�4Ei2�J��L�Q ��N38f2(b4�m���E��@���3�#4&D2�����LQ�6D�x�y\g�����k������k��ɨ� ��!�!!��� �%3&<�o��[�j�� ���px&����ry&Y�wD�a��<�/�<�� �                   �<�o!!!�/� �%�3�o ��p�x�o��r�yoYw��&�nEi`F�n�J<�/�<�=�/�=�Q6���N��݁q֠3�X?�,8X?�4qdq!.�/�q�!3�lD�aE�`F��t����Q���DiP�� ��3�2_b�n:'2O׀�;'2�J� �                                 ��݁8ք��/o%3&_&32&/�"//b�o� ��'2�J�/��4Di���E���/�� n%2&_&{	&��6	c56b!5⠽�2�Jā�8Ki/�& �ꁜʞ p3/&_	&?D.�??b	/t�ǫ�x�y�m���%3&<liY�wD�a��<�/ቭ<8f4oYw�E`�F��<�/�֪            �=��:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&��:�b;�h�:&�;&���:�b;�h�:&�;&���:�b;�h�:&�;&�l����=�K ���� 	8��U��x�� � ���/Z�� [	� �����y�!"⨖�y!. �/�y� y&��y�k� ����r�y<d�x�!⠪�xyf<�KxfFy�k �3.&t�o��� >�_&{	&��6	c56b!5���.��֪t�O)��>���Kɚ�)��t�/�u�� �3B'_C'�p�$

8�4҅�� 3B{rC�}p$ 

�8�-4�- ������~/6]~'�-g�h��L�����ڎ9րC�4/�hM��ssd�ɨ/~'�����7vi����������ɡ���ێШ��B�?���9�nC04/&ssd�ɨM�������� �                                                                         ���bD��槦"��b��b�!.� /�� �䍀� ��F.
�!�� /�����         �����6�����6��  㾿k A���'��0�c��%0��bJ��
.���d�邾�r���"�d�ꂾ�r��d� �    0A p                           ��݁<�xyf$q&%3&�:&�;&[�Yw�Da�<�/�<��X�?* 8Xi?4&X?� 3Diaq�����x�y%b3oYw�E`�F��<�/�<��U���x 8�y�4�k                                                                                       ��݁<�yxf%3&�:&�;&[�Yw�Da�<�/����%�qXi?* 8Xi?4&X?� 3Ei`F�q�J����B��88b���풶ڄ�!8⨸�� ����

c��b

�
����(� � �  ��"
��@/���� ����*� /������c�o��c�&!�뀮� �?�������              �Oc���C�8��@S�  P� �A1����Oc�	�� 0�0 ����O�c��H�4T` � A	7��A�6��A�5��O�c��0�0�C�00�C��0�0 ��� ����Oc�NXQ�@D	�R1�D  4(4Aq����A4����Oc���P�0�0�A�>00� ����      Oc�NQ�� N�TP U  � 40&0( 90b��8.7Ai79	:A�9>	?A�6B	CA�5F	GA�8K	LA�0M	NO�c�`00 �`00�:�00�:�00�cB��0L00�0 ����� ����7Ai7_	`O�c0�0�M`!� 5 � O	cҕT`!R� � /z77c7/b|--c-�k ���r��/.�8�5�/( 6Ai5�	�A�6�	�A�7�	�A�-�	�A�9�	�A�8�	�A�/�	�O�c�`00 �`00���00���00���00�cB��0L00�0 ����� ��4�(94.8.7Ai7�	�A�9�	�A�t�	�O�c�C�00� �`00 �R���D�0�0 ����� �