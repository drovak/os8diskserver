����� �C : �B f -���������                                                                                                                                                                                                                                                                                                                                                           �������7�&��)��/������bb�������� ����)����J�?����*��?�����r��s ����0�����0������&� ?�����c(�����&� ��О馞頞��f� ���C(�� @/ـ���B(��X')���FGÀ� �@� �����������R����p�2c�����  0�
���`�����/�֮�l�?����*���!.b�" n	& 
�
	7�J����F��&�B&�(/�?����r�~&�C����!㨸�!.b��s�&�2c!���&��k   ������:�7W)Vɗ �_�S������� �����l�6�6�6C!�.c�������f/��"�b�&"��b�b���(���(/���!���,����/���餀��颠����0����< ���&��!���d�J���&�/����k�"H��� �          ��	�a���	0#O� ��?������o �i��S���,�� ���r n&�	&�&�É�4	t�����/�����s��s��s��/����v��0�(?�����)�(�����?!.�?��C�����)�>������8����� ���Y���� �� �1Yw��� ��h�H Y�@������������_���������F����� D��!.��b���F.���&�(?�����c����9�)� ���7���q.��/����&��6@./o!NJ.

���&����� �   �ǲ�&�����i���\ �   �ײ�&�/������� ���꡸HYW��Wx>�whB1��X�������� � �)
  ��� ����&�"b�� �
��+D�.c���� 


�� ������������������b���˽(� ���b&!������"�����* ��������� ���8 ����᠎���� ����ᴁ�!����;+�X��H���
s��p>�w��`?������c�&��D��4�JN
��	&	
&�/�&
	7�J� ���b��&��/�����|��'��'��'��'�� ��ⷷv� � �� ����ר/��/�٦�{���X��
�������)��?ꃼ� �    �����������k�'��� �F����vɢ��p �p�������� � ��( ��,!�������)��"������� � ���������� ���t� ���7�����b��s��b��s��b��s��b�|� ���7�����r��r��r�|� �      �����u�&Ɂ<ꉜ�(/����b���/�ɤ����� F��f%���o솀��9�������X������ @�ހ  ��&��) ���"�����)�J� � �	�����������{�
��*������/��"b��

d
(?��
1�����)
�9�������t�����������+�P���)�h�   ��֣ � � ��                        F�@R��HH�V� �ɇ��`���o ��>�����0�����S����0�����) ��������"������������y���E���� �          �	��0�����������Ø� ��(?��c������9��`>�?�/������v� �      W�x���P�O���Z x@1�Ywh�`��'����` 솀��� ���c(������ ������+�����b���!�⠺��2�&�	&�&	7D�������7��� �� ��l)��  0��� ������ � ��@?ڀ��"�b!�@��d�É���Dܯ�����J��� �   WA̑            ɇhY����0�1����������� ������0��&��<����t��D�����c��ǉ�Á�ǉ�ĸ�D��J��,��r��|��ɻ�"�����'��'��� ��  ���� ��� ���Ɓ���(�J�����F���� `� >��b�8p� ?��"�����'��J��� �� ��         > nb����8� DL#� � �L#� � ���DM��C L �D@`XaS%@��XA �R���DDN�N E	���e `R���DDN��TUR�C�@IR���ETN"��TUR�C�@I�8�l3ɂNB� R���C	��TXVCm�P	$�@;R���CT� E��S�$N�! S`	 �A��C��18CU�T N%E �L�S�`���N� N$ 	Q��@�e6 �  �TUR�C�@I�T�D�E3 �8�N2 E���PE1 ��� R�3L�	T`��PL�TS@ғGN"LRC!�T��ŖDD@ON5 �ShTT �UE3� �            