����@ � �+'=>*'*79!>+'=>*?: *2'<: *''>/% ;$9!>+: 8*8: 99; <+1*'=>'<; 9*.   y<77%6(z   ?2<(*?                                                                                                                                                                                                �����2�����̨�� 7�����2(����/�����~��x����� ���ɀ ��� �� ���É����������'��'����:��̀`Sr�݀��0�H��A�3�N�G`����d� Љ��Y��A qO�3�T                            ��������%�V]y� @!#�0%f%/&{�D��z����n0/&`0�%#D���� ��(�b
b���Z�& 
 ŪJ��� @�6�b�N�/�F��&�F.�� ��(��b�b

bb�ن&Z�& 
� `�6�' ��tׁ�� �/�i	a>�/�	�a���	a>�/��� � �~ �� � �0�o���b�n��&q.8/�H�&/&{�bb!���&&��a.�/��������a.�/��������&������j&&��/`i��bba���'��r���'�����n&����������66��J� �   ��ݟh� ��(Ͽ̦��'�J.�������t��"�F���bH����&��&���J>

�̓�̈́� ��� ��'��D�����t��'��0J
���b������ ���R@����$��t�]�                                                       � �����?  �$ O� ��� �      ��1l�;\>��"    �     �           �          ��O�        `        �  q�         � ���^�B���  @0 R� �����$d�" ��(����� s��@ ��M��8
me���1b��$�o� �gh2ꀠ��`?��8�?������3����k ���f~�&� b}�`����$����t|�����F�����⺀�D�@.�/�@�(��@n/�"�򺳊 @�/�@�/{iz (��!�⠺���!�⠺���!�⠺����� � ��F.������r��/��最�  y�/�|��خ xb�n��u���}�f���� <<w)}�v()<} v()�u�ts�r�q:p ;)b���o:�F�n')m~��t����r�w���lk bji�h#&#68fgu�f��e��d2�e�u ���/�خc|�~c9�c9�c9/c)2c)ur�26/6�7�7~75�J9e�gK2�Jb��{�!�����a��&��6`g��� Cg� F� �C ��)�/�_�c(��^�/�]�(]�(ݘ�&�&�I���J���G_&��^�(��3�"(���(/��� �����Jv &�+��x��n 6��+�(��+d^2(���(/������� ��
&
(?�(�_�z�����b(ai(k� kw	�?�������2�ހ���? ��/����1��!��\�1�B^(/�[�'��������� � 1Ĩ/������1�Z1&�1���1�b'1��Z�1�h1�J�!.1Yb4f(?�'�4X"���ŷ*8( �"�!�����')!�(���� ��b��f����C(��@/ـ���B(��W')���W"'ӛ�t� ['d�'� X�Yb]b�t��� "!\i����!����7o���50ba7☀�7/&�2&�V�VV�0a./�/�{��)�)�)v()�(�a.//&��2�J[()75D�\�7@.*�ɏ�_��       Z&F.�.qW(��ȫ )(�����;J.W�(:�W()�(�/UV)�(_�?�7�V���7� V�[()7�k@.T�� ih�%bl#%!>##$Ȓ�#%'i��iS�%#b!%����#%'R�l ���ih�%%c�k�Ӑ�� �� �� �� �� �/@!.$�jF�������f`i�0�0/d$�J �       � �� �� �� ֱ �� �� Ϡ �� �� �� �� �� Š  /��xQ()[()0a./�/���{)�* ��*����(����s(����s��������zP�)�������Á���������������'��Á�������7���|�<V��
��t���t�����|�������'! �����6��C��b�(�o������ �
��$���ނ��d��� �N �-��K"�W�& �
�!�"���?��k�)�����'�lx�wk�)��b�������/����Pr�����/�Pr�ȟ�����{��#BA�DAJ6N�RG5�Dԏ�CQ��Á������kà����'��D��J�����|���*���O�΢��w�a�$���|��8�0�_ ����dB� !��(�?0B��!@�������}R��_�����Ȁ��(?��'��Á�������Á������!>��/�����r��r��y� � �	7��J��� ����z���"�*�.�1/b08/ ��%
��NB��A��CF���̳����b��b��k���8�O��� ���h��/��&!��^����d�*   ~,�(/��kr����$t	c%� �)����ɥ��%� }�V�  Q��(?Ǡ/�Ͳ~��-"-�b��/�����"���N4&�v�ͣh4q ���� ��O����F.O���7�J.
�O���r��d��J~�)�Ê��&��B��ry�/4 @� � �
    k��b��b�@n�u�N�*u��� �M�/|��� ���y����J���� ��|������J� ��fZ��_�صvw�|؞3�h�y�(��v!.�f|������� �(�3�|���3�a�c��  �� L"K�� B� �}����J��w����� � )��� ���?�I�''�'l������~ /�ӂ�*�   �
� �       a��b��&�K"F�H���&�P.��/�� � ����G �   �G+ԃ&�%L�G5S  F(/������|���u� �"(����/�f�À�r8�7bJu��a�c��+(/��+|i�|�ur�5d�a�o�bk!k ���t�b��bj�gd�2b�� �"(����/�ؾ�|�2�J&b�bbb�j!.�/�a�d����w����w� pp (��n')�H��T�.�\��@ ,8f5�bc�,�/� ��J.����|,� M"(���(/���@ ���/�f��E������Z�/�a�c��  � /� /� /�(/��Ⱦ�e����K#b� ���/�#�DD�%b#%D ��#&|E��#�b�#&##6#e��|��*C^�/��|i�a�c�� �khPoH���4#� w�3���U1�d2��/�a�p2��5�)�/�a�s�� �y�/�u� �/�,����.bc.�cf���d2��ਵ�(/�.ui�,�a,&�خr�.66k (��!�k������8&?�A'��~�&.} ���az�.n ���l &#6# � .V �a�i��k �Dbckw��D�~��ז" b�J.(����H(���H.(���⨟����5�/���5f�A���� ��!#�#$���!.��wn�b �� �� /� /(��C�(���(/��(����R�)b�����J����#6�#+��B��z �(�2����"d!)b�\�[�&������@�� ���t���v`�v��U �>�@��4V���)r��Vz�(����)�)!.�/���(�!��[�(�� �
�b�b#~b
w#�J�k i	(��h�&a.��6��bk�j����&_c9_�sRi�D��T��_�r��&��{ur� .&�jJ)����&�J��' ��&~a.h�6��hj9h�2�� 0S�O�Cȏ(0k� 00p.@�/����c�c`i� �H��B@����(��n��(w��V��� �   (���@/��"�)���� �����/"�N�/�F��	&�F.���o� � /�	�	c	c	c�lĀ���)���� �                                    ��! � ~ �U; ���%��� ���)�:f;+f"?f>f3f_�rmi~&~j)�t�)b(�����_�?�]�(]�(B�s�����\y>�(?�(\��P��
�lkH0
=r

w���T���|*�   �c�(O�V��v�'�������   �ڥ��'&�(&k�'��j )�/��P.TI���彠����E�S����7RK�"�&�p2���|u�,c)c)c)�c)r��Z����66,6 �" ��|�� ����9%��9���� �k (����b�nbb��bwh�#�b#%6�!.#(?���%!>��/�%���J�w)S�&#!>��?������ᠮ#0����#�##s�%&�%'�!.%�"� ���b��f��&C&~�*       S�F�W���"�uir ���/���u��|+�!��+�+b��+�"��� �"(����/�� +�+_g|����"�uif�����d��/�a�p�� a	c ���|�� /��	r	r	r	�|� �#�n&�"���#'���k�G+  �@.��/��K E	�f���� � �"@������%
�F������	�D� �󽲠���k w������z
�
���i � �
�k w����bkD�k !�敾&��8��4O���8��4OJ
��

�󦊽�O�����    ��)R����X��Yr�4v��&��Á(�*� ���kw���6�&�C0 H�Z
��d��6��F�����([�(� �l���q�n����vr��uur�)(/��8�7b�]r(��w)}��#&#-"-#b'�}'	#�!.b@���#�J�#��縲r�&_{�/�����r�!�&���"5f�!�)�/� ���|ɚ���X��Yb
�j��J���� �
�~|i �/�\�)�� �u �F�/� ����� ���K��� � � v*&��p��" #�#�H�##c��ˉ�Á
ΐV���|�����Ⱥ�L�����Ⱥ�C�(�J����"��� ����Á�������'��'������{  ��'��� ���/�*�k�/�~�*�d�*�/�J�()Q()�1�� �k2&~()2�J����LR � X� 0Œ EB$�T�Y ��J!��/�@���8��������*�
��.����|��<FV�������'��Á~������'��Á������u�����㳠����'��D��J��́*�q�����)�����'��'��'Էr��w��'��r��r��{�aI�⋪0�B4�P8���=�n���� �6�O��WmLg�!�"9� F�PF �
Bl�.I�.\�J��£����� �M �  Q���Q� #�錣 ���ˡo6�.墼��e�	��SǓ� �S ���S
��)�S���(�猃'��煃�9����Z��ŀ���e����e�	��ü��E��=� ��7�tW��x�⇐�˱zX�� �   �`��+���� %�ޠ !�o� $� &꼡  �ޠ "唨  ټ� �%�  �P� QӼ� P�%� ��u� �%� Hͼ� �%� (�%� @�P� �9�  �� ��� 
��� �ޠ �ޠ 	�J� 
��� �ޠ ��ޠ ��J� ��o� �ޠ ���� ��� cޠ `o� \�� Sޠ S�� >�� ;��  P�  � �%� A��� ��ސ ��� �J� ��� �ސ �o� ��  P�  
`  \�  \� \ސ No� 4� ސ �� ��%�  |�� |%�  {�� @{%� �xހ �x%� !sހ �pހ ]S� 3��    �  � ���b�Nb��lǁ<��tǦD�ɢ���'�*���H0(���*�  ��*�   �
��y�~"�V���'�H>!��6�d��'��'��'�ɳC��ɳH��˥�������GU�NU��U��UA�|�@�!&�/{i�� a�`i/&D�� ��
.

�l'	�} '� ���u��'�xR�k������� pa9&Ɗ��=6�h� ���Á�τ)� �� �&~')�J���s�@-�T���(�e�����7��D��J�����s���Ļrźy�R�pl"I�/���W��  %��U �%                                                                               �	���!���?��#�@&@@6@!.��s��������n*&����cF�����/�����&���wt����d'�0��&&z0��~����t����7�7�76���/���T��{���[6=����j}�� ]5�� �       ����� �E�� ���ں
��_                                                                                                                                                                                                