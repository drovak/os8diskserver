����   � @ 	  	 	  	 	         >(. 	2: =8 99 >(*4: 99:<2?: 2*)98/#<;?)   : >(/;                                                                                                                                                                                                       y�2 R               ��� � î "3?"��!!�  �                                                                  b� +$                              �70 �                  �90��ǩ2 � �����������������Ië���)�����������K ����� .��d��J��d� �    ��@ �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ޓ�(��@����)��J   ���� ���&��'� �       �@ �?p?�/=� !�  !�� ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}to�nm�{|� i_@IQe���r��������i�����g���ˀ��������d������� � � ���������y�����y��� �����Q�!@�?>="��"��"��������6��H��h� �   ��)��9��� ��?�>��� ������������������TN"�  �	���/�����)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP���3>"  M�À��"�"=?"�  F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�f���� � 5R�� @         �� �����"� �� � �� ��� �����A������l���Ήl����������������)��"�����"�����"�����"��������������������'����� �ρl�'��6ς,� �   �� �LD  �� �C� Q�� 茀������            �   K	��� �   ��B ��
 =B�kX�    @�       ���̀!��'�\� ��i ̀שo��l
�` �d��ty� Y� I�5�+��@�P�        � $  h  ����?U� ����� �����C�X �                               �	'   ��
�Ĭ��o � ��� �������{��n�nQ"��b�;��<'�='��2��89&� ��Y��c�:"($�"���c�+$��� �����=!.�r:()'��+'� �� YB:"(��!Ӛ+��!����:()�!� �� Gn":()@�&*��v���nc&$"����+c�$"� �� � ���� �� �pq�� ƥ������  ��	�h6b��� 	��h6b���� ��h�n+���+� � �\]f\h&])A�]�O\\B���]x"��� �,�6O"\�n]]bh\b\���\\&�\���]�/�]��� B��?�!��\]f\h&]){�{����]"]o\\B���]x"��� �`���� pR\&]�^�_�`�J�Ia&^h&])��`h&_)��a�J\�J �� U �Y�n+o�c]f�\6]�#^^c���]D.()$"����+]�\�J ����+�]�c\]b�^6^�?�<�oc&]D.D"(*�$"����+o�c$i"���+�o�)$���]�\�J ������N���X�5�8S ��"�H� ���Y����6
"\�n+؞<c&�D�:()\*)��$"�����+�h"(��خc$i"���:�(c�$"����\�J ��*� � M�hiH�*h&H��� ;��M�h&X���h&X��� I��U��R�\KbM�h\bP3:4'39{�*�h\bP	{�*K)���\�J �[�*����p.  �R\&L)Eh&\P 3:r43s����h\bP	��*L)���\�J ���*K):4'3Mrh&���+��hi��*K) ���*L):4'3Mrhi��*+�"hi��*L) ���*K):4'3Mrh&��+��h&��K�� Ғ��  0��6��'��'��K  c$�� 7rq�R\&K)\P 3:r4Mrh3c$��\��R�\ih&\P $��K����\���  ��R�\Lb\�P3:4'Eh&39H�:\�JR\&h�\P H��L����\��� %��R�\Kb��:4'�M�h\bP533sn�����h\bP5n��K����\��� I��� 0          ���� 0�H>R\&L)�:�4�~Eh&\P 53'39��:��h\bP5���L����\��� ���R�\Lb\�P53�~:4'�M�h3cΓ�\��R�\i��h\bP5Γ�L����\��� ���R�\Kb\�P53�~:4'�E�h3c���\��R�\i�h�\P 5)��:K)���\�J ���:n:"^Ui�R�\Mbh�nP)/�Jv�&\; J�^�-7�-\P �|�]�mE(/�]��E�f\b;Jh&7j&\P i'i���\�J ���:U��R\&hPb_��v��cf\; J^��7��\�P�|]&�(��f�\; Jh�7j&\P i�j]�J'ؚ\�J �2�JH\&�+�M�h\bO	��Kh&\O ���w���~+b�c�k�(A�	�D,#����\�K �`�LH\&�+�K)Mh&\O H)��Jh&\O H)��Jw�&�+�pb&qc&,#����\�J ���LR\&L)�:�4\rP53�~Mh&39��J\�JR\&K)\P 3:r4Mrh3c���\��R�\i��h\bP5���L����\��R�\ih&\P ���K����\��� ����� bTR\&L)�\�P3:4'Eh&39I�Z\�JR\&K)�:�4\rP53�~Eh&39I�Z\�JR\&h�\P I��L����\��R�\i�h�\P 5)I�ZK)���\�J � �ZU��+�h����n:"E()�E�c6b*؞-�-�-'��$�"� L����+�7))n:"M()*؞-�-�<-)'���+��	�c7b)n�:"(*�'��$"� �i�ZU���+�K)3:r4:rnM"h7bjXi�c�7�-h�-3�=���E� ��3�Zh4E4H>���3x2����E�f3cio ���Z� �� �D@�:IbZYfK):4'3Mrhi��Z��:4'Mh&�� ��
c&v�&f")����+��hi��ZK) �� P���U��\bn:"h�bB�z7bjXi�y�\�i7b�h��\���ݙ�ffbE�/�خcfb	��v���jy�j���u�&K)���\�OhhB;��\�x�/�� ��U����y\f]b:n"hXi7))h()\*)'Ԛ$E����\�Jh]D]�/�\�x�/��K)�u�v��o �E�jU���y�\]f:n"hXi7))h()\*)'��$E����\�Jh]D]�/�\�x�/���K)�u�v�o �t�jG`&^�_�_h&^)��jK)���`�J �� `U��I`&O�Ha&\�]�^�_�K)_:"4^r3]rh\b��_�Eh&^)��j]h&\)��j_h&^)��jK)���a�J`�J ���j� ������ f�U�s
�{VI`&\�]�K)]:"4\r3y)�z]E"h\b)���)�z]h&\))�zK)���`�J � �z�`&�PR_i^n]]bh^bL��_��]�h^bL��K����`��� *� U	���y\f]:bnh&X7�)h�(\�*'��$�E�/�\��h�]]B���\x"����K���u/v�&�� O������~)}� �bO !d⠌�e!.c�/��K�}�U�
\&�`&�_�\^&K�*_H.�R�
\"^LbH�]afaO 3^rDH�337��:4'4E2h3c���a�=a&]�J_�J�d��_�\^&�_�H��R
"\^&H]&a^bDH�e�oh�aO e)��zd�/KK"���a�?a&]�Jd_d�\�	\&`�J �� p�2�n���+�k & �R�&��d�अ��� �\i�� �]]bAD(]�H*	'��+$����\A D()\H *'��+�$������9��8�9�i���������E�����}��2�/�/�>�������+Y�Z�k�  ������ �V[&�-�-���-[����
-)iib��� 	�� @3�3�3r��� E`8b_�f�:�H�+�_�J�8b_�i:H.�����_�J��_`d���8_&�:�H颈��_��� ����� 2	/�2/�p��8�c�2i/u���"��b�)�)�����&�)�!.�@.�����8�C����J8�/�8�!8���h� ��= ��&�= D:�� N��?�溰� �       q4<H�� �`8b_�g�:�H�+�_�J�8r_�i:H.���v���j_�J�:�H����c]�b>�&L)�:24]r34sEh&39TҚ֓h]bT��L����:�H�`����8_&�:�H�Ȉ��_��� ���� � D(h�()�c�$'��خc$iE�/��D�F����� �mmb!c����ž ����� ������ ��\�Y�\�\\b@:�� �]��� �^��^���\G F�/�_�\G M�/�\�h]bԙ�Ѫ\A 4\rh]b3_r��])�Қ_�/�h���^�њ�^�� ������ �(R���f������������� ״'������ �   kkbjkb������� �D@�:�nZYfK):4'3Mrhi8��C:"(*�$����:4'Mh&8� ��
c&v�&f")����+�h&8��K�� � 	�� ����� ���6�B���ڢ�´���r�r��r��r���    �XR���f'���¤⽤∯��K �����f�f�+���~�/²   W	�{6�����������d����2i2��A��o�/i2�/����0��Dﴀ�/ꛀ�/�b�1c�0����bD����/�d1)e0)�����&�&N�&�@/�D���b��D�/i�0������������+��+����D����D�J�8   W�e   ������������ �-
�-g�gl&l�+ �V[&�-�-���-[����
-)hhb� ��7�Sbrgr�J� �s�n7&Tr&s's .rt�B��{�i
������+h��(	�+� �h"(� h��h�+���   	�����$I.��)ڞ-,�&%�2��+T�� ��n:()hD"n()�*)'��� ������� ��y�z6�hB�n:()7))�*)���c�$E����u�$z�{t�*f	 ����h�GF���y�jv�* A c7k&hA !k㨻�hA �k�k!>i�/�i��֮Sr&kkC!c���c .crd�k�B!.k�?�B��خcyb����y�vz'�c�kl6��K�NĀҀԀN�̀���D��   �V[&�-�-�-�[�J�
�-e�V[&�-�-�[�J�
�-O�d�k [[.
A��9[A �9� ���������� �  ��b��bA���d������ ����ɵF�I0(��@�
�

���J(��@��)��N����@�� p���&!��"���� ii�-���� ���� ���6��B�:bn()�+� �ύc΍dh; n:"D()�*)̚�c�R�&$E����Fc&fC"���h"(ڞcXi$'���F�/����Ѥ�̪�c�$E����h� (c�$���vB΍{t�*    ��An��"F���
.��&�/�x������b��&��'�>"�n��sH��� ����� @             � ��X�{6 � �����������;Y�/�Z�{��+����K8 �c7bkhbA!k�?�h�A�
kkC!i⨶�i�*k�NTr&k!>c�/�k�c .crd�T�rcfk�?�k�r�Jk!>B�/�B��خcyb����y�vz'�c�kl6��K h � h��������T(}�E�d�8N��N���MM� 闙��'��&� 6 �0� 7��E�������!  ����zw��m�jZب�U��U�V-ffdD@DBEDH�DTSG�S%�RA��D�MN ��A�RA��� 0	����DG�S%�RA��D	�T�`R��D�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C S��P5   E ���� Gb��v:b=�� .99b�b����9�bD:��/�#נn��tةJ98&����@�  ��E�����6��Q�&�/���À�P � E������}dؔ�Q�&Ϻ�������b}�k��� @�  � PP��@̓0� 4                                                                                                                                                                                                