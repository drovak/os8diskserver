���� � A8  
 > 5>���������                                                                                                                                                                                                                                                                                                                                                         	� �@ٔ�MA    !� 6_� ˀ     �                                  � �               +  ����� S�O�^�UB��� R@� � ����dB� ��(�?��s�@: ��M��8m�e��a��$���g2�� ��  ��/�>3�2�������
 �	�������/����/����/����/����/����/���7� H7��H/�����y����/����/��j"F���e���#.B-�i���-����e���!�⠺��������F.������r��/��會� bx" �!���/?A04�;8�V�� � �0�~)�&~��}�!|���{Á��/   � �"#f$%f&'f(zi�(/������z�������/����	&�&z�����	'�J��K2oft� �"����d�|��d��d��d/�d2�dt�q�2c/c�s�s�5t�9�e�h2��c��z�!.�/�/�b����nso�!�Zf����� y	�b
�b	cb��/�
��J!.
�?������ �*O��yb	�l�<(��b

�
��	r�	�O����<���D�*���/��f f!�j � (���� ��+ z�����z������e�/z~��"���z��(���(/���(����/��~ܚ�?����Zv��? A�!� ��	F	(?�&�!�ʀ�� "��������!�h-D�.�-�he�K ��	F	(?�~��1���1�b'1��[�1�h1�J�!.1Zb4f(?�'�4Y"���ŷ*8( �"�!�����')!�(����N� �b��f� ���C(�� @/ـ���B(��X')��� X"'ӛ�t�O\�'e�'� Y�Zb^b�t��� ��/��������+�3&�6&�!>�76�F.�7"h��J
�
!&5 �  p�6����6466C�6��J
4�

�6�3�J�F.&�����       �[�&�F.���.pX(ٔ�ȫ    )(�����:X"(������W��`����7W)V��7 /W\�(7� ��UT3 ���f ���b��l{(?����������࢙�b��l���@eݚ��{ǁ��,�b��r��r	�l	(?�/&	06	16	(?�2&��¾�l��<��   ⾢|�r+�b�b*�l����D �͊,��� @�΢5�k������;@Vxw������ �� Š  /��xR()\ "���/�#��� �c� �6f�b3�c��r��r��{ ���x��hb����t�.�ଫ'��D�������;       +��,��  `�����b��d���w�K�ȓ�����;����װ�� �� �� �� ��  � �� �� �� �� ��  � �� Ġ �� ҍ �  �� �� �� �� � � ���"� $�T#  ��� �� �� �� �� č �  �� �� �� Р �� �� ��  � �� �� �  �� �� Ю �� �� �� �� �� �� �� �� �� �� �� Ӻ �� �� �� Р �� �� �� �� ҍ �� �� �� �� �� �� �� �� �  ��  �  � �� Ϡ �� �� �� �  �� �� �� �� �� ̍ �  # � ����>�3�/�����r��r��y� � �	7��J��� ����z���"�*�.�1/b0   ��%
��NB��A��C "΀� �/ �/ ��" �BT < ur��h��/�ⲲP��_"���e�*��~,�(/��lr����$t	c%� �)����ɥ��%� }�V�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                