���  $ �,/*,+$  =.  
$(  Z % 	   %: .7=79<*.**77<7=	2/
/79*7<
/7<7>88= *08=*08?*0'?*.-     %?  .6	%	      	 	                                                                                                                                                                                                  
    �MA�#;�!�� �                   8 ? ���� �� �� � >�����ˊ ����������� �p6 !,	S!�� �  P ������������������: ��9� f.?`[ ` 8    &!f�"d�k�'�dp�: #    bm�a����  0��M� ���c��b

�
�葒(� �  (��@/����1� ����*0 /������&!̧������ ��  7�d��d���s!!��� ΀��!>6�/��!-⠵�/d(�� ����7b	c!	��� ?�������� bx�/�|��خ wb�n��u(����}��� B�� Q�A �:B��A3�8�1 �
B��A3�8�0��JB�� 	Q��T�`�3 B	� ��:� @�*
�)�&. ��b*��&.���"ˬ+   ���    ��&�	� ���b

�
��� ��&�. ���&� ��&�. ���&B �   � �0a�h �    � �� Cg� �
�=�����w��� ����B� H���AB� ����2�B3R � ����B� H���AB� � X� ����B� H���AB� A��H��@ � ��-B� ���A)B ��C�M% � ��-B� ���A)B �	IS� 8�"�BiR��DS`0c� ��0X������2�ހ���?Bc��B��Q �U@B	c��BN�T�/ C	7.8�g�-b!8�(���#b!8�Ȍ�$ .8�?�8�
)��8�����/����}6 }���}�iB���T@� �C9��� ��  �
ɀ�9Ґ��  �
ѿ�9Ґ��  �
ـ�9Ӑ�� �  �⫀9i�� �� �� �  j��[ `O\�'e�'� Y��Zb^bduUcUv6�n&.!.�?�#�!��;�& .�?;�(�a�c/<��J�J(/""f@.1$ ����>�3"!�+&�(�@�O=������ .b,&A)B��1 �A�B��0��C�E���C݃c �C9��� �  :컀nc7W)V��7 /W\�(7���@U��7�����q"��fȸ(�J5&����� �b���и(��(۸(�J��(�(���S��h�J�b������w��&��� 
1E&DE���� 
2E&DE����H$8 L1P1 �T 0      [� $� _� $�$ �$$�f 8 j 1 � �"����b�k�q.A � 0�H>�����|B�� E�TB���3�C�׶t"������Ԗ����������w�]I���ZI����FJ"�\��V�WZiJ�/xW���ZiJ�/xZ�K�/xZ�L�/xX�WZiM�/xW����.ZiN�/x��X�WZiO�/xW��Z�P�/xZ�Q�/xZ�J�/x��Y�WZiJ�/xW��Z�R�/x���� [F�&&__b?`��q��-�����2�W�m���W�J���w���������w]�FFbK�/�����w������_�怎怎����!������]�(������`�栎��_�N_?)`�mw��J������u"������]R���� � ������w�  �-B� ���A)B ��TR` ���&��_fu"�_�?`���w2�W�m���W�J�b�GK������wH�!_�y�ZZ�Z����w]�a�!�������w�HHb�z�Ha)��w���������w*�ab�]*�/{��w�GU������wH�!`�y�������w��_�_?)`�mw��Ju"������]R����"�	 }�T��&���t"����������m]K ����$�����/����ۀ @   �&&�tb�-2W&������W�J����W��]�K�/�W��/y�&�J����]�R�/�����i�Ի:  ��b}�b ����J�}'��K   r `}!>�/�}�ܠ���j �)|������ ���_�ص�[6�t��-����]�R�/�u��-2W&������W�JK&7	&����W��]�K�/�W�	t���B�` A�B� K7b		cAB�� ��J:��u"������]R���t"�2�W�m����W�ϖ�C9��� �� �  :��u"�2�W�m���W�J����]�R�/�t��-������E&y%M�H5S ������w�������w�������w]�FFb� �������w�������w�������w�]FF�+ FT�/x��J�/x��  ccbb!Dc�bb&cJ.

�ccbb!Dc�b] b�k �������H��]�� ���6�0����6��[��C��zd P}n
 d� �ɔbFCq�T�*�\��@BŔ �TT� ���@SC����m�ߔ��������r"��b����������@��H��Ȱ����� �   BŔ?T �	B)�TB��8T��5`�3N��`	�3���LD!��� Ec ������m�����ڀ�ᒳC_�/��|i�b�c�� �k�h�PH�� �4�#�� �y3��[6 2�/�b�p2��5�)�/�b�s�� �x�/�t� �/�,����.bd.�dg���e2��ਵ�(/�.ti�,�b,&�خq�.66l (��!�l������8&=�A'��~�&.} ���bz�.o ���m &#6#\� .W �b�i��k���Dbclv��D�~��ז                                                                                                                                                                                                