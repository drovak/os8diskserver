����   �                                                                                                                                             
     
     
     
     
     
     
                                                                                                                                                                                                                          ��X  ��  � `�        	                                                                                                                                                ��b��/����<����9�����b�@/���J��/�̢�D�y�9�6��"@����������� D���"���˓��(/�����������9��9��t��                                                       $d�'���P���/� �ݓ�&�/���F� �������F�� �	 ���B��/����������:��&�b���� ��b���F.� ������D��i  �� �	��B��/���I��� ������̀���RI�2(����/�⭃��                      �� '�� "/�5/� ���C��m�� ���� ���������f��&��"����=����� ����D�������&��"��j��2�����2�����-��K                                                                                         `�e ���  C�0 ���C��}��0���� ���������b��f��&��#�����=����� ����D�ɤ����&��2��z�O�������r��b��f����/�����-��2�Ԁ �                                                            ��eq ��� � �3� �����ڀ ���6��C��d��6��C��d��6� @��4  तt �䗁�� �    ����!�죠?�������!>��à����J��� ���̀ ������̀�����                                                                                 ������b

c(��!�⨒�
�J�/
�6 ���/����H�)�������

c(�����
��i �

�J0���(/���(���/���                                                                               K�7��
@0 ��E�Ow`US�HV`TA�1���(�EO�4���_ ���r��I�t݀�`6�Rgǁ4`�6r�{��u %V`��3`��AA  �R QV`!��C8`�%�E ��O6`�U�8��6E�t�(�`6 � �I6��;� ���`Sb̓TA_ ��I�c����RFI�c�Ѓn�k��p�`6N �Eg��A�	�8�4T_ �?%���E�UC�H`��8R�XE!�ԶR`vGI ��7�R �T�3]���	�]Ρ�l1�]T�� K�8]�	 eX�o7  ��O`e��S��RQЃ` `�KAR���D��� Xo�#]�� ;V` �AA��4K �D@ ҵT_! �]�S� AR���@ P�KA��L�'��X�8A��p�5�8S`VR�� @MR`� RQ��D ��EÃ��# RQ��D � �E��C�qT` �EgUSA �VAu����7��XU�RA��D � LNb�DS�R�� @S�(��3 �PPR0@� A�@� Dt B��@�@@� @�@�@�@� @�``$�j#j$��$��$   ��ª�c��F������'��2�������� �� }��                                                                                                                   ���&�����c���������%�o�D>Ș�&�������_�������0�&�,��|�'��'���b�f�)���!.�b		c(���/�	��	�k!.�H/"b������)'�J�)���&� �  �          � � A�`f�Y�8������ ���n�)�)�{������������r�h�������������)�)������)�/����rc��&���k�)�����󛃅�� ��%��������   (?��ڠ�&� �                      �����Pޤ �e��
 �/���������&���k� � ^����  � ���d��6��C��d��7��D��J� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���&��,��恿��J(��öj���J
�
n

 �.�����l� >��b�|p� ?��"�����'ÒJ���Ã,��� ����8- 0                                                                                           ���&��6��B��f��4 ���.�(����� (������� ����(/��(��(���(����"H���)�����&���Ük�������                                                                                 
  � �?�@� ����l�!,����&,��������,�(/������̛����(����/�������                                                                                                                        ����}���                                                                                                                                                                                                