����  �?% $<$>%%%%%%%%	%%%%%%
#��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                   
 � �MA�� ���L �    8@ ��     � ��������PH��(�       �Id�3�� ��̸ֲ�ΤG� ���� $�(,�04�8<�@E�JO�TX�\`�g ��EK�QW�]�� \�U�"�&*�.2�6:�@u�xa                              -P�- ��z�l�n:[�ŉڠB�[ǝ���l�nI[�ɕ�W���l�oi)[˝�o�i��jo�� �[͝���lobi��jo�p[)ϯ�lii�j�op�� [�ѹ�i��jo�[ӝ�o�iU�jo�[՝�U��j�o[	���oi)���i�j�� �[ٝ߀�ij�[۝蠮i[���ڠi�j[�����X���� (;A�U�l�nij�o[	��U��l�n;��=��?��A��@��ij�op[㝘�Y��S����k �  ��b	�b
!b�c�
c�
coob p� �	(?���� ��J� ��&�	&��&!�&�6�&��D�
& �&
�6
o6o .p�k ������	(?������૊�ݔ �       �   ���� �    S	����o�;��C[����W��Ǩ���o=)�D�[睒٪X��zl����o�?��F[����S�Y��Tǘ���oA)�H�[띰٪ǀ��o�@��G��[흻٪Z��� �ob�p& q&�&ln&o .oob�lp���ln&pq��o��Ǥ� ���b���� /��@� �P? ?`��؇��� � S	'n&lTi;c�hC�[��liAc�]H�[��Aa�](�)[)��W��l�i���))A �](�!)�[���������8�A� ]	H[�����X����l�i���I); �]C�[������'�l�i���X) ]	D[�����Y��l�����g�; �]C�[���������s�= �]D�[�����Zߚ�����" T	�(�)�'=)u?)� ��6��Co�d�p6�CpTy� �o�J� �Se� o&llbnld�o���n;)]C�[����W��l&Tc�hG�[	��#o&p�fpq&��&p�JoO��� ��b����&pl&Oq�nqb=��?.�`]�D[� ����l&�n&F[����T�l�n=?�.@�]F�[	��X����    S	c�����'=)o)&u?)]H�[����W������T�'=)oA)u?)a]�)[)��X������㙂��h�6����b����/��㨠��D������>�*�!&�!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0�H> S	�O�n=)p?).`�q�l�l��6q�' �� ��'/�H[���W���� wo&b��f�!.��b�!.� n��b�o �����������&�n&� p�d�o����"� `��/�p�!u�������b�����J��&獢�l���/�듢� N q�<�� ��� ���3      
��(��H��� S	l&E��[����E��[��W��_�l&?)G[���G�[��l�V?�G[���X�������)߾1���9߾I���Q�ʾ����� �ɾ&�?�� ���� 9&��9�/�!��"�9�k ��;i  ��mi;�  ���6� �� �4�i�4��� 2{��{Ɯ2�J�����2 S	��� lTL� �[����ek�AL� [��ꄠ�lTi;e�h]�AL� [���T�?���eIk � ��L �[!���T`�L �[#��T�fL� [�%��Ta�bc�L �['���lTihG�[	)��leikA�hG�[	+��Th�TG�[	-��W��lTiE�[/��� �R��"  ���&#UTTc�dE�[	1��T?�@A�E�[3��T�hE�[	5��Tf�E�[7��X�꣸� �lTiE�[9����l&)Ti'=)u?) A�b]�E�[;�����Ɋ lTG�[	=����lTi =�^8�.`�>G�[	?���T�>^�8.	` =G�[	A��Y��逵�^B���]&s~�v����~v������U��T��� lTE�[	C���lTi'=)u?) A�b]�ek�AE�[	E���lTi�=�^8�.`�>e�kE�[	G��lTi�=�^8�.`�>E�[	I��Zś��6� ��fE� ������p �B�
� �2�J������� ����p� �2�J � � !.�/�� o�g� S	lTiK �[K��Ҩg�oTi  [�M���W��Ҩf�oTiek�A � [�O���҈i�o-Tiek�A � �[Q���X���e��<�T�  [S����i��H�T�  [�U���Y���� ��d�o6��Cp�dp7p�7� �o�J�v�JK�LJ�MP�QN�L �)�nA'�=u�?b�]e�kA�� �KG S	0���fl�h��o�Ui^ ��[�W���W��l�Ue�kA�^ ��[�Y��l�Ue�kA�^@��[�[��X��lUi�^� �[]����lUi�^���[_��Y��S�� ��6��Co�d�p6�Cp�{ o�ҫ � � �֠�� �@�  � @o �
2�K �ut�yz�xv�������� ����3 S	leikA�NL� �[a��éf�oeykA�  L �[c��ĩ�l�=�ND�[e��W����l�n=c�ND�[g��éf�o9Ty�;�e � C�[i��ĩX���R�aHgǞ� X� ���y ��2�����y՚e�y~�z�2�J����yy�~z��z��2�����z������?�. �� S	l�h[k����W��l&�[�m���X��'�l�n)TiA'�=u�?b�]'�=��A]�D[�o��)&l�b�Ti'=)�*�[yq��Y��� ��n�)nbp�h� �n�J�O��� �n)&n�"pnb�D!p�p�h� ��O���D�����nd������ ��&nn�"b��k T	pA)'=)u?)b]�E�� �    ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ����� ������K ��ʴ� ������K ��� ��� ��� ��� �� �x b��&��mmcm�c�mb�\i���V��x�+x  ����u�u&"�|��'��'��'/|��{���1s��}�9��o�1��o�/࠮~|f�}��"b��b��b�f~�&�.��d�D�����3)�1y�����c��i����������줮�������B3�4�71��5��1��}�n{2k � �e�       � � ��r�~            ��y1i����=�,�;�W<�� ��}b����s� �6��|&��.A�?O�%	 D����, ��!.�Pn��ݦ�� D!���"��isK�,� �y�i=�,�;W� S	6ߒޠ���i,�sK� �	([� �� �� � ̻��$��EEbFGb<<�b<)F�JZ<)DO�E�*� �!���� .! �&��� �DhF�� �&�&��h�	 ��O�D��摷����/3��4s�1yǿ�s��v�� 8������&�6�� � ��1顾� ������8)��"����(?�@��梠����j��Dʀ��$"����%"�����C��b� `���������� ��?�'�i������x �� ��7'��6��?����V��|�/����|�d�1��5���(}2k ����������&� ���sR��3��R9��r3�4�7�!B�"b��b��b�Xn�o�͠�����b������6�����X���d��J��'1˞� ����� ����   � �   � Ѐ����R���Ok$6�# ������ &2����� l��� �m�(� n��� �Cؘכ D	�C�� �FؘC�; G	�Ƅ� �EؘͯK H	؄�� �x�(�� ��I��v� �ʉ��y� � ��& ��c��c� ���K ���6��0��7��C����t�3)�4c��t��'��B��t�p�    : � ��t��q?�rns�l� 6/!��"��{�����(/2��(2���/2��t�/tv��v� m&\���s�z⠬�r +r, e����   �}�t6��Cvtbv�/�l�?F�[������ �1����o�o8)o$"���o%"���o !�w6i�b�\�f_�	jb�
ne�rh�vk�zn��q� �# ml!.m�/���\�{y�/�������\�s��r7�r���V���K+�e����������5��6iy��P� 4�7��nz��w�CCb8 �����J���c���C/���������/� ��{�f��{ir���x�x�xd�/�4����������� �z�w��<����67�<����= "]O"�62 ���&��&��&��D��6��7��J� ���⣧b��b��d��C��c��t���� �    '                     6�̤�̀�̌���������g�q Є���� ������ ������ ������ �������� �� 5N���@1�N�� 5�N ��`1��	�8 ���6��CR����8��J � (����b��/�6������/"�8)� � ? ��� �!Ϭ{����{�b&�Τ � ��8)��� �8)�8)8���  ��bRʘ��b��� �� ��b�����+      0���R2C � ��A3�8N`!�R1�� �DM�P��HG1L*�����D 0	   ��� ��z��� �{�/�!���{lAO�Ԍk � � � �+ � �K � �k � �� � �� � �� � �� ��&� � ��� @)��� �����&�@)�����K   ���?����K Q	  �� �h��;]�� �F�������� �?� � � #� 4� F� g� p� ����� �      �;�=?�A@�<>�    C	�D��F��H��G��C��D��F��H��a�bc�_`�de�fa�bc�d��Č����������������� �A� B0 C0 D0 E� F� G� H� I� J� Kp L� M� N� O� P� ����$��$��$��$��0H� �� ��0��0�� H� (� H� (%�!5�%�!8A%�B%��5��! �1 �1 �1 �1 2 |||�||||	2|
2|2|2|2|2|2|2~2~2|2|2|2|2~12|22|A2BC�LD�LE�F����\�\����Â �"(�"H��7�3.#�8x`1ϔ� C�TR� c\�I��C1p-�mc  �S  ��L�C ��D��ЈS�    � �� R1��D � �T�H�8I�PR�Fc& �Na EO3��O-��  �          �                                                                                                     +5D��D��D��D�EUHJUPRU��U��U��U��U��UԆW��w��w��w��w�.xJL�������:;�=?�@<�>C�DF�GH�EB�IM�LK�PN�J���������ę�ʙ����H�49 ;B DF ါ         ((�  pp�pp�pp�p(�$  >                                                                                                                                                                                                