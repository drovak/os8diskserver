����  @	.   	? (/)   $   $ $ $ &       #;?  5=���������                                                                                                                                                                                                                                                                                                       ��LT�0v&xş��C ���G �   �� �� ������E�?D0   �&���(ˁp�   ���8 �t�C ���0���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s�
��� �v���؇?����� ��)��)���b����������)������.�i�����  ����� ����r�b
�b��y����T���
�~�b�f�� �� �
�&(?�	�6�&	�0!����J¾��D��耾� ?�!��� 
.

��� ��o��3�� �À 4[�C3�/��D�����4��4�&�&���2���J�/��"�������)�������i����&�	&����b	�i��)𥉉�����
&�	&	(?��	6(?��
'
'���
�r� Z�&�	&����Z�/���k� ��i��bi ��Xp���� ��$��(�B"߃I8��E�p5�����	&H?��6	�	H?�!��/�	�!⠊������)���/������&�	&	�?�	����		&H?�	�	7�	���)�Õ�����������r��r�b�bt����b	�j�
�	(?�
�	6�&�H?�!��/����@��b���� �/&���� �S	��($�2�����YB���q>��/�����(��
t����������i�"�������󛍍���� 	  ���	  ���������/�� �����/��� ��0���c��0H�����	r�	 �	�{�+��D. b ��?� � ��������U �CJB����5�?5۞P6P cbȴ�H.����/������"���J.�n	�~F.	'���H.���H.bJ��	� F��*�	� ��bg�J� ��n&��c���&��c���!>h?���&&���H��� �67'�(����H�s �=m)<�&�� 3��� �Ϡ��	&
&
q>	0?����ھ�{&H?������D��tCt�J ��c�������6�C�����)����?������i�2��C����� �>����&�c���(�8���k 
.���(� ����雰 ���3����5ɞS� ���"��"��* ��&��  � ���D�J� ��
'�
'��K��(��(� � @���(��� ��߰��� ��(��� ��ʺՈ�+ ����/��� � �b b�  b����(�J� �&!�׀��˺��� ���(��(� ���(�����3��Ɋ� � ����� �?�� T��� �߀d��6��Cڀd�>܀d�H.�
n޲h��ʔ���(�����ۍm�F��&�ۂH!��@/�!���ރ-֕� �!�⠲�܅-�� �����-��"��҂��ʀ���K ������,��/���͏���K         � ����dB� !��(�?0B��!@�������}R�}�� � ����E��_Ќ2LS��$�RFE�$�TS�����T�5��; �� ���2	�4� @ŔsR��E�� ���H�8RQ(o�� 8�tə���XM�P�0Js`��8	� �Cp�%`���T�D	��ON5.Q��wTL 	ϋ��Ҡ;�@��V`��Vn! S�"�@R�A #�B3R υu��MW�F;Մ3D�����Np� 5��TS�" �R���>NTO�# �0 ���2�N.�R�	�F��`1SaQ��w��T��� ���2���`1��  �Rp��3��� ���2N(Se`R0A��8�H��D�MAS���'Ѕt��S�`FN�U��AD(��5 ���E��4`�e��AD(�)1�� �S���'R���>L ���m6�TR�S	�4�AԏDE.a��wC�DKTC QЅt��S��C� ��WqF;Մ3 �W��M D�0� H��3 �T@`�T "SRW�S�? X��s_ ׉tE[��0`Vl!��	2 �YTR��; ����DA����T@��RQ����_Ϋ` �  ������  ��  ��+|i�|�ur�5d�a�o�bk!k ���t�b��bj�gd�2b�� �"(����/�ؾ�|�2�J&b�bbb�j!.�/�a�d����w����w� pp (��n')�H��T�.�\��@                                                                                                                                                                                                