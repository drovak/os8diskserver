����@  6 *$">6f   2	?2>=<9
9
;:= *998882	726=/98
<(*"8*:288/
:)28 )
+ 8< 
1> *:
)*"28!;> . 54. &1 g4;$?/ :?6. ?? >6A                                                                                                                                                                                                � �      �=�                              ��            ��3E�0��      0C� ��� ��7��@� ���ЍZtW�����0 ?VD�k3��� �:�� ���(�/TPA���V�^A��� ����?���
r�o  �&�䶻�n�6��6��7/~b�g�/�}�b �� ��@�␑��"�|� �f�(���(/�{� �� ��B��b���骈�� /��/�����z)�"���y�J�*'�J�"�����b������y��"���~r�k�
������ z (��~z ~<&eww����3�/� �� f �� f!c�@.x&��wB�!bD!� . o�����!�*��D� ��/v�Wv; ���4�ui�ģJ
�
����4��� t (��|t |z)�ò�y�� � ��s0����K�ċ �r�&�� �q��pb�{ �l� �@�o��
.n��/ぼ:�vk��Ư�tl�i �� �O�y�e��lm�����/�����!l�~c�� a."�/�!�a#☫�k� b"!b#�lq1&j�1�&a."(��H��!��lq�&`.�/{�"��h�/��� l'!�'l&��Ot�Ѣo�&�J� ���i2����J�o"�d�ޢo�&��hۛ�g� fh"�#�k�� �&� !!��)6s'k��q�&@�&e��qbh�?s��/��&���{"��n&���{"��j'���.�d!��c�EO3�H��T�5L�TD �T�	�3σ΃� �ћ��b��/��@��@��(��@��@������Bt��&��� �E���'0t���������!�c��hbF��0�hbt�00&�&C(O�0����6�G�v��� �4P�?��k��m��=�g6�{��{과�������;��;R�   �&F>�2���ya��b�h�҈�H�y�� t(|'`0(X�7D� �     �  �� �  �   v �  �c@._/^�" ���a���� �B�o��'(3(3((3&$373<3ES3�i�(��p&�J�o"��j|�*���.�.n �֢�����B��]J
��] F����b����b(��s(π����\b��x�* 	�8M�P��Oyy�y �DT̓A�3��� 0 D SK :B AS IC .W S  ��E�	0  ��/�d�Ѩ/��`�~�i������Ҩ��$��%b��h��������b�[b��lZ�    ��-&�,&��/�$�(��(%b)&b*'b+�k��/((/�$�)%&*&&+'&���r��m)� � $%&f�'&�&w&�қF���қ7D�ҫX��Z�	�
���dg�   �Q$� ���t��/ fqb�vY&�&ț&X�����_�(��&������   o���ț&n H
�
�r�]t�Kd,���� ��Oʴ��dYY&�&��d'��K� �M����8�8G   .����n�b��bco6'��t�Jo�"�d�ԫ�M�m@P� ���LG��|�'�W�V&U&(?����~&�J-bЁnT���-b�Z�   ���'��'��lZ	�d��d���|`�-�,Z�$  ������!.-�/�Т-[b�-b�Z�  �ǲ,�lZ	�dg�   f&&�q�1ci(/�p�a �(�����OeS���e�a>!(/�����0h�S�ё�� �I4Dt�y�������j�&��7����nWr�c�WuW��/g��a���!��u�g/�����g�z��    ? O^ /��/��� (��^ /��/��� �                                                                         \zx�z�P 3��a�����j��1��rb!�����(��!����b�d(?�������C闊C(��颊��~&� .��j������~���b�b��b ����!����D��J�&�(?�����J�Ԛ�К~rc(��z��y�~&�������Jb�g ���t��"���� �      ��*���Ae6S +��         s��@.{@/�@/��/����В��/�Т�����)��"�����K��&�(/�����s��(/��� ��J�������� ����@>�(/�@��@/��/�Ј��z�� o�|��o��Л\z)~&!.�/��z�܅�D@��w����w� pp ������3����@��^`��� �	��(��\�$� �t�"�������l,'V��É�(')'*'+'��6��� $ �
�������d-���&�{0�v{ !�&������DM��C   ~&�&^2�����Ht�����] ��7��B�]���t� �4 ��t� � PH���	7�&�����O�W� � �����s���̢�Yb�b�di�(/���,i��
 �
�dI���좞c]@J
�c]J
��d�4s�(��_�+b�g��bc(c)c*c+gk����������T�d�a�&-�,Z�   Z	��(/ݚF����dv�� �+d��������Z�	��~����柎b� �a���!��b��g� fqb��y�2������j���q��rb1b�s����I�j����q�'��D����r����F�����'���� ��!r��y��r�s���Ԛ �'!�'vK ��s�(���(/��J ���/�d��������O�3��o�nZl�ka� �+�Q�� �a����!�␌���)��b���|�z|�t��&��fw�&�0&�&@��0D�ꤜ���&@���.�/�O�D.��&��"��d�ꢠb�� ���n��b���bn� ���/���'4z���� j	0�i(/]p"�de��6���                      0   [k���`�ԃՃ� 0o�#R���C��S�m �� �      DS K: BA SI C. WS  �
��ÁZ���������|�����&�������w��w�&��t�f�y	(?�Ц�����   ������|ȁ����X	 �
�.�ǁ����d����+\�� �   ��������P� �������� ���<b(��]F��
&�&
.�����&t ��/���'
7
7�J�NFBMRAMKYJNJ[LA[GS[PO�N�D;C DH�LP�T ������� �D�� �� ��������FN� P3XSe@�?��P.TI���彠����E�S����0\�6��"�� ���<���0JJ��%�@/���F����ÁZ���s�H
(���j����l� >��b�8p� ?��"�����'�J��!��⠀���'��� �?�%���J�w)S�&#!>��?������ᠮ#0����#�##s�%&�%'�!.%�"�S���b��f��&C&Y�N�o�: �����