����  @?8 < <?< <>?<>?>8 < <?< <:  =< <:  < <;= =8 << <; ? ><< <; > ?<< <; 0 >8!><< <; ? ?8!?<< <: = *4:		< *2$: 
3)'40: 	8	> )'		0&0!*?0                                                                                                                                                                                                 
     � � ���L �    ��       0 @` ��  � �"  4 �f Ϗ�������������������U�  � ��������7  ? ����?�j���`
`寵 2�K���Z֩A=�.��� �(���. /�(��+� �(� � ���g�d��( /�(��&� �(���$ /�(��"� �(���  /�(��� �(��� /�(��� �(��� /�(��� �(���<H/��.H/��<�@���.@/��= . ��?� (�?�  ���> .(�> . ��=�  ��� ���=� ���G.� ���@���@�.����@����@�.������+��� o � /�� o�  ����&!>� /�:��&�'�!.� /��U PP� ��!.� /�T�a� ��!.� /�^��	1G                             ��b����&!>��/��!�⠈��� ��b�z���>�
����  �������̀@ �����d��2����ӊ����P.��/�٨�!���0��O�٨����J�ъ���ǀ������6� ���J�
>

�堮��c��@��b���� /��@� �P? ?`��؇��� ��.��@������@������=� ��@����  ���@ �(���@ �(���<."  ���;+"  ���:("  ���9&"  ���8$"  ���7""  ���5 "  ���4"  ���3"  ���2"  ���1"  ���0"  ���@.�./ ��@�@+" ���@A�(/ ��@�B&" ���@C�$/ ��@�Q"" ���@D� / ��@�E" ���@F�/ ��@�G" ���@0�/ ��@�=" ���@�.." ���@<�++" � ��@�;("( . ���@:�&&" � ��@�9$"$ . ���@8�""" � ��@�7 "  . ���@5�" � ��@�4" . ���@3�" � ��@�2" . ���@1�" ���@�"2 . ���@�3" � ��@�"4 . ���@�5" � ��@�!"7 . ���@ �#8" � ��@�"%"9 . ���@$�':" � ��@�&*"; . ���@(�,<" � ��@�+@" ���@=�/ ��@�"F" � ��@�"E" � ��@�"DH" � ��@�"/ . ���@!�!C"K . ���@#�#B"L . ���@%�%6" � ��@�''"@N" � ��@�**".O" � ��@�,,"P . ���@@�@<" � ��@�==" . ���@����@� ���@����@�.��@�=� � ��@��<� (���@�..; .(���@+�:� (���@�(.9 .(���@&�8� (���@�$.7 .(���@"�5� (���@� .4 .(���@�3� (���@�.2 .(���@�1� (���@�.0 .(���@�=� (���@�
.��@�
. ��@�
.��@��
���@�=
.  ���@�
.; .(���@.�
:� (���@�+
.9 .(���@(�
8� (���@�&
.7 .(���@$�
5� (���@�"
.4 .(���@ �
3� (���@�
.2 .(���@�
1� (����
0� (���@�
.(���@�
<� (���@�.. ���@�� ��@�����@�=.  ���@+�<� (���@�(.; . ��@�&.: .(���@$�9� (���@�".8 .(���@ �7� (���@�.5 .(���@�4� (���@�.3 .(���@�2� (���@�.1 .(���@�0� (���@�+.��@�. ��@�.��@�����@�=.  ���@.�0� (���@�+.(���@(�<� (���@�&.; .(���@$�:� (���@�".9 .(���@ �8� (���@�.7 .(���@�5� (���@�.4 .(���@�3� (���@�.2 .(���@�1� (���@� � � ��@��(���@Q�Q� � ��@�L.L . ���T.T . ���U.U . ���@R�R� � ��@�S.S . ���@ ��� ���?�.  ���@ �`� �@� �� � ���@ �� �@�P�@�P�P���� ����� ��0� ���?�. � ��?�p?� � ���p � ���?�. � ��>�� � ���?�.0 . ��0�A � ���?�.0 . ���!� ��?�� ���a � ���?�. ���>�. ���0. � ��0� � ���?�.0 . ���0Q. � ��0�Q � ���?�.0 . ���?�.0 . ���1. � ���1 � ���?�.���?�. ���q. � ���q � ���?�. ����<� � ����0 . ����;� � ����1 . ��� H.4 . ��� D.7 . ��� J.3 . ��� F.8 . ����� ��������� ���� ���<� � ���0 . ���;� � ���1 . ���>�.< . ���>�.0 . ���>�.; . ���>�.1 . ���X� ���X� ���T� ���T� ���Z� ���Z� ���V
� ���V
� ���>�.� ��?��� ���?�.� ��>��� ���?�.� ��>��� ���?�.
� ��>��
� ���=!.0 . ���0!.1 . ���G!.2 . ���F!.3 . ���E!.4 . ���D!.5 . ���Q!.7 . ���C!.8 . ���B!.9 . ���A!.: . ���@!.; . ���.!.< . ���!.(����� �����!� �����@�����!� ����P�����!� ���� ���� ���� � ����7� � ���� ����� ��)�3-� � ��3�/ . ����� ���� ��`���`��<�`(����� ���� ���<�/ ��>� ���?�/ ���P ���P��.�P��.�P���� ���� ���.�/ ���.�/ ���0��0���&0/(�� �0���� ����� ��$�� ��+� ���p��<�p��.�p��<�p(����� ��<��� ��.��� ��<�� ��������</��</��<�/ ���.�/ ������� ���h ���<h/��.h/(���� ��<��� ��.�� ���>�/ ���� ���<X/��<X/(��.�X@���<�/ ���<�/ ��.�� ���.8/��.8/��8���.� ���.�/ ���� ���<x/��<x/��x���.�x���<�/ ���<�/ ��.�� ���� ����/̀�>�/  ���.D/ � ��$� � ��� � ��<��(� � ��� � ��L� � ��&�,�  ����  ���<�/ � ���� ��� � ���� ��� A� � ���A � ���>/?A/  ��� �� �A� ��� �� �A� ���� � �A � ��>�?��?�  �A�? . ��?�>��>�  �A�> . �� �Q ���  ��� �Q � �� ���>/?Q/? . ��>�  ���?/>Q/> . ��?�  ��� �� �� ��� �� � �� ���?/>�/> . �� ���= �� ��==  � ��?�> ��>�? ��0�>!>/ ��?�?!?/ ���@���W�WWb �����W&g0��W�W�W�/gX�WVb&!̿"�gǠ���͠�ӭ�����Ǯ����ˠ���ō�������Ԡ���°�����ή�̍�����������������������                  ��┓b��d��������&������� �    ��� n��,������C	���MN �̀3`��R1`6N O�3�TN� PT0B# � �U� @��A5: ���D�E3: ���@	DA�0��0,�� � @` �� 5N���@1�N�� 5�N ��`1��P�@��                                                                                                                                                                                                