���� �= --19 :   	     ( -8/ 	  	 2.1       )%( 	 	   -8 
                                                                                                                                                                                                �+&@ٔ�MA    ���                                                                       ��� t�W��?���� ?V������������� 2�K���Z֩A�?����� ���� � ? 
 0 ���� `"��  �����������?�!f�(?�~�.�c(��~��?���}�?���������&.�,� �
�/&��&�,� �
�$&!�/�����f�.���   �
�0&�.�i�ך.�,�&  ق��־����|/�����l��  ��?䁬�u�|) �&0��.��ҩ�?������ %��n{���z� �Iz�y=&�x�+$i�� �� N�#&���#&b��/��!#㠪��J��Ⱦ���)���#w9BF�w��#"#�j#w9#+D�x�+#b��/�"������w+�����������z��Iz�z��{)�"�����Kt�c�%\�� �AP�@3*��(��#֞/:3 2����24�k�2����2
.ۄ�4| F�42b�v4�2�

�ۄ�2.�4���2
.

��2���4���2.��2�
�ۄ�4v F4�2.|�4�(2
.
��2�ۈ� =��/��K ��&� �u3�����{3���/v3"t"{=�=�/���{s�{r�{y�=�k؇>�<�E  �9�d�7&9
>

�9��9�� �q(�8�8�"(����/�8�p�78"{��s{)r�*7!.�7&� �H���**�+ ����0���g�&��<&�H�x�o<<*r

�o�7B��/����/��� ����ۺJ ��� b ��l�Ub!�l!t=��!�z���;� � �`� ����"&�%&���n�<��� �h��� ���f�,�   ��K !���z$��mÁ�ɉlÁw�(��k��z�8�Kz@����������� �� 88
.

��8�� q (��pq p{)� �}�8&�c�'���8(�c�)�� ���b

�
���� q � /��/������� ������.��  ����2�H�	7�J� ���w9�J� ����J�k �P� �A	��J� ��&�	&x&� ��/�z� B�z��K z	I�L��<(��:zi6:B�z��K 11
.u��1�oF��&�7�7z1�1v ;�l��<v!;�/�;";�cwJ
;���)�����&�F����32D��C�� �
t{6�t{)� �65f6q.5�8?�!��665�$� ��!¨����:�(?�~�;;c�l� ��(?���6�6n(?� &�����m(?�!�"%f!lCw(�k����mH>!"�m�H%�mH>!m�� �+�"���� �-�b,-b�--bv�t{),�J�Ժ���   ���� �� �ֈO����?��A�4��8Tz e����N �z�AC�H� q�8�Li@�� 8��w��2��wGm��w=8�^{Cq@������R�$�L�ބC� ��s�z�AC�Hx�C��Tp`���p	����AM�RQ��C��` � ��Rp�4��w�RAe��AC�	H�Gp`��sހ�T@D`�g� ��N�B^R^ ^CY�N�RL^PG�TP�Ԟ�1C���J�j+�/��������� �      ~��A�i~�	��� �L6�~	�� �                                                                                 V�X�ߟ��