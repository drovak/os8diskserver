��� L B    �? �=��b�r�RS�(�!�r�b(���J!p���k�8�   � �W �      �{�����2B)��ʉp�2B)��ʉ'��`�������B9�ρ �.B)� ˉ ��&�&�	&(?���	R9-(�¢�/b?�����	�J���?���J�7 �d�� ��/                                                                                                                                                                                                �������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ  �
��D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �      �����}���v	P�n�_��F ��&J.
�����ȳ��������R.�i���b!�⨫�Ȁ����}��  0����&W ��&�@�|"���J"��&��ԉ|����/�C��J��b(���}Ɉ � ���k��hB�?������Ի �?�"���V�"�����'�N��PTB 0��� ����� �� R�` VV�!�ڠ/�F����ڶ��r��x|b�i�(��m�������(��m(/�@��|��i�����m(/��������z�� �"�b� �F.��+�(/���H��bV�������m /���ڨ/��� ����� ��c�(�������F�߮�!������?8��W��2d�pD�F�&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{   �(?��B6� � �gWq���� g�t��D����/���}�� $����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ���������  @��      bH�
��bmF��B@���Pn����� ���O��O��������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�޴�����2X��(?�
�

��������������o��R1��D��� N E��D� �@C� ����	��T P�ل�MA	O���� 0���/a�   ����b	�n	t����w�d�V���T� � � �? ����]���aOY����&7�B!!⠌�!�6]Z9Xc��c'���b��&��7��b��/����naa7�!.�`bc�t��!&`!>S"���O0�����b!a�@��a�xM>]]s��/�O�MT�a'�!.cc7]rG�* a�`b�f�?��`!>&�2��d��          � � ����6��6���H  �� >������cJ���t��7��C?�F�0�F'��0��c_���t�6��0�c{(����m"�m�m�&�m"�d��&�lሐ  0���k �&�9 O��J���`/���������n��&� �    �?���b��kG�t�WF��&�������Dd#pD