����A @?=&? 7! ���������                                                                                                                                                                                                                                                                                                                                                                 D�@���� ?��@�      �s` ��� �� �� �� �� �� �� ��  ���ߟ� �+�Z! �!�
FZ� .�� 0D����.+            �� P � |��b8� �,D�
��U��U �
8)9m'm��� 0 �P       � �G���/ �}��   � �K� �8M&JHd&=b?UrVfrv}v7)�7)rtf��"�Kf+6�@5����K�t�t�h�� DI&+ט�0br�(t�rtb r�@b�srb�b�I�(�4 bŀ�� �� �� �� �� �� �� �� �� ֣ � � D���4cH��!D����#��c��k׀N�׶}KBFK��♢���"��$��Q��"٧$��B#3��" �D��TAo�nBa␪�"8)mo�r�j*r��r�r2)LJd�LÁP� r�nQbGfY;�a��� @y"�b�D"H��`/�����D Ȱ������ G�ڦ�q"�ǁq��F��q nG�k ��Fd艬�<bbb

�
��F�b @.(���ݪ\�$�	"z(/��(��X�+n�3��fI3
,(�/mo����m*� �Y�cA,搐C�Qb{�/b��   Tr�nsb�rb2L��L�OOcLOr�N�s�Jo�/n�boo&��n.(b�r ns8bMJd�m� r���}�/bo�!s�rrB!o��b�r2)L n�L�cPbO�l F�rn&r1I7�����im�D"���s�JƯ��A	ON)s3Km;�$"<@�.&�@�DAirnDoB7Q�Gf+;�"<�� D.�(��7)D�+ !@b�KKbo��b�R�*�IÁ �IKd�I�������t�rbF�b�Ef@r������&�E�@r�r .@���E��8)�FD�m���( D���;��pDBMڛM)p#b��M��uȟ�$��J����p)"@��pbMp��ګ.&�>?'Q&G+b,�3�33 &!�ʀ�� �����+��"ާ&H�I!9sbfe"ee"� P�˺������L��� z�(j��H�ZM&4!�M��w�<�m�ZM&�&�u��M���J!��m!��H�����]�0rr(�!E�/m'0&rtf}Jf�S��E��Ԯn9bmm{��A�� �� �� �� ��  � �� �� �� �� �nr(/nr&r�r�2� F�1;�v3E�!t�ȭ�x .t�/bE�2s�x�2r�t2)t�lsK6rs7tr7Kt'�m��!"I�1"!Q�G�/H�/,ҹ'bE�lQEsG�J��� G� �Ecq�,�	���E�zH�.B �FYi�/�D�IFd"D<iIC+r!.t�/br�Etbx:k������ù19�!����D��Cc9�� ۯ0��W�/b��rhbV�rc�k�[+'�� ��i)7)�հ r!�so"�b��n�o�KDf}�K�  <��q /QrLPrQQrLdQ&G�l�߸!��w �����o��H����Wv�m&9m'wc&w�'8M&H]B0�t������U�܉�w�<�b�o�/���m�k�)����|w� ����DDb(���ȿ^U��vc����n� �
� �߳�ZM&�ȿ_ܹm�6c�&m�&�����#H����s��cx�lxH�  �_���`���	����c('�8ך��>���n�����m&�m'�c&� �   ����� ̍ �                                �� �� ��U{�S� @x!l���8x�8����	�k�lb�n�+�kl��!��9m'm���b�k�Bv~rWb����߲�k$n�JtnTk�J@Q�{�/�Q�!��t&�9��r�b�-Q&onf�Rǁmˋ�à����6�<� a�,��{��s	�p��8��8��8��8m��� �� �� Hk�/�����b�b8J�+;��@��J���D��zn.nb!���g��/��n2)L�f�L���c��ln!.o�/�� nF1i��b�/�n������ª��/������䷊��JF�/� �& F���������/�o���no��K ���j �c(��!��褰         u��7��vw� ��&F�F��2(��Ҡ/�F�!���2��EEc(���E�b�*�P�Q!.P/bF�� η&7F�J��QQbLb�L�� �3  b@nb!.��/�b"���MJd4!�Mm� ���ڀ��t:+���x�&!���8#�8
�8x��8)�i)j���*	!��m�i�e�  ����ȿ���5�N%L�G�U�&�&��&�Éǖ�Jf����'r�l���   �HB���D�"�����K+�2���� ���L��<�����7���7)�7)��*�M� /��/��"��gd�2b�� �"(����/�ؾ�|�2�J&b�bbb�j!.�/�a�d����w����w� pp d� ���p�Ј� �e�� �����ŉ���� ���'��0�����ŉ�����/�����,�|�.����6��9  ۙ���� �o�(�����������/������)߁���f�	��ぜ��?|�l��/�&��d������I	���	���	��c���  o��W�������U� Z��K� w�3���U1��  ��?��!����&ğ&� ����¨��������&Ơ/Ӂ��O����F.����7�J.
�����r��džJ��)����â��d��'�O� �   � �   ���щl��0��&�?ǂ�b �ǌl��&��É����ǃ,� ��l�����'��� �o ���}��  ������~��ז  ����b��l�(?���������� ���r��i��K��0�����0��z؛��Z �����bP�␽���̍ �� ��騷�&��K ���l�?������)��������������!�����2(����(������ ����� еF.������F���G@�?E  (�U�  �����B�k    ������J�/����&�6�(/���� ���0 ��Z
��d�6��F�@.�/�o�zN

���&��̞ �� �ν���&�� D�� �bӼb��j��O�خ���᪏�&��0J
�
.
��戣����C��(����$������U�������f��� �                                                                                                                                                                                                   