����  @            
       
`                " /"?!#!/#?  " " " %"'"/ '"' /"/ 7"7 ? 7"7 ?"?#!##!#!#!#!!#!%#'!/                                                                                                                                                                                                  @ٔ�MA�� ���L ��� �� �� �� �� ����D5�D��3]�� 1 7� h�Pw��gP���C"4�  ��<$                             )? Q� �� �� ��     H������������������������ ���v���? ���?���R��` 5�4�6�7�8� ��� ����� ���� ����� ���� ��ߣ�K ��� ��� ���� �ߵ�K ����R�Il��������������N)���& ��I��M)�_����� u (��|u |)�ظ� �� �(?�r�� , �d�Cl���YC�BAf��A��B���'Y�CE&Fi��E�JF�JU����������������������&P�Ě ��ʚ ����"�i���� ��ޚ� �AP�CrR�	1G                       � 1"��#&M)��C�B]bABd�A�����ە������[������o� ��[� ���$&M)!�C�B]bABd�A���̚���C���������&�� ���Z ��_���� /��@� �P? ?`��؇���J� �H�HZ  ��H�[ ��H\  ��H�] �� �H�HZ  ��H�[ ��H\  ��H�](��� ��HHbZ ��H[  ��H�\(��H]  ���� �H�HZ (��H�[ ��H\  ��H�] ���D� b ��l�Ub!�l!t=��!�z�<"�i;)�f��H/�K�dC&*<&<=&h/'a�'��7J-BGeb;%k�J�KdBC)b<<b=jb/ar��s�er;.bG%kȇ�q�9�/���{z$�8��)�7��6)q��5&����9�/�8�I�� & 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� 7��3��dC&�J�K�oȒ�'<&f/'+G&_�*(<&g/',G&`�'��7e;&<=&=>&e:&��������YC�BAf��A��B���'Y�]�!�l �>����h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0��3��� ?]� ��C�DDd� �@?b!@�0�?!.>�?0>�9:����CE&Fi��E�JF�JU��\���� �l �l�������Y�;�����D�D�J=�N%Ի�����d��6� �   �ۢ�݂��d͊���  ��� ���d�� �v �J
�
��(��H�� ��S�W����@��J� 7�K /8���?@����� 	�;RR)��:R"��>S��?R��@R�� �&!̷"���� >!G���<>&�����5��  6�U��AP^�U��BP^�U��AP^�U��BP^�U��DP^����!�����!����B ��� ��.��
.

�
����   OX�� H �洹&��&��@��/�O����X"����d��J������� �   ���@���e�:i��:�Jʚ�� ���4c��b

�
����(� � Q (�� Q� ��ޛ Q�l@/�Y�V�ޛ �U)T)������ �LD!����΃`�G��D�8 �U��1	ES�����`�LD!���D@R�8A�'����LD!��A��1	��T�>�_T` �GD�� 5�S`ǁ4`N2�TP?U U��� �LD!����΃`�GD�# �T? Pl�_R ���	�U��H��AM	�R1�D�����DD�� 5�A��@�H�`1�G���� ��@� X�@� X� � X�@K� X�@K��_��4��?� X�  ��_A�tBS��	�U��H��AM	�R1�D����N�A S�T��C����A� ��:�������D�:�M5TO�8S�8��DDS�HS.�����E�UC�H�8��DA� ��:�������D�:�M5TO��; !��E�UC�H�8��DA� �R(�.i(��D�(E�A	5�n:�C��A� �R(�.n`*�8STãMTPO�#S�ԃ���DAS��TS�.�_Z,)�+�[b,��+��\,)�+�]b,����@	�0T`     @ �   $ I���F$m�����"�#M�3�4Q�DUU��UYf�g]�w� xa���e���(i���,���0�q���4�u��8y���<}��A��� E���S`�w�BLT@&XR�� S�"��3��@��T�` M Ք3��X�D1׋M��h6-���C��ă �01 23 45 67 89 :; <= >?  ! "# $% &' () *+ ,- ./              	 
   01 23 45 67 89 :; <= >? 5@
�    ?                                �   � �                     @A BC DE FG H� JK LM NO  ! "# $% &' (� *+ ,- ./     �         � 
   @A BC DE FG H� JK LM NO �{����dB�LlxW�J�A��W�U��p����9�����?_ۘ���ip��v��v�7ޑ<;$2�|��~ �       @�/��G׈o�������%����'��/��7��?7��?��D��N��ǈOψV׈^߈W_��e��o��g���w����w����
�����6��wψ                                                                                                                                                                                                                                                                        