���   �?;?,#���������                                                                                                                                                                                                                                                                                                                                                                       ����c�����DрJ{�,����{���|  �����r��r�b�r(������c�J
���@.�/�Ӥ�������"�rJ��� �&�7J.
���&�7�7���{�   /c�s�s�5t�9�e�h2��c��z�!.��� ·��p�:�F�����	?$	�D���V��f�&�&����/�����bt���'�J�"����"����)/����)�&�&�9�J��/�����)��)�������� �  �  �����CV (A�`   �  �  �  �  � �� �@1          �����b(bi(l�4�l�AMC�@3`?=���w���?V  �  � ΃`   ��S    �@A   �R    �� P   � F    ���S   I�  P �� 0   �S    LVN   LQ� P R%N �RNQ ��E� 0�FE� ���SE�I�NQ ��5N Ņ�`6	��`F ���`F ���` Ʉ`fŅE�`6G�`&N�T`�#� A12�34�56�78�9p�qr�st�uv�wx�y�̱�̳�̵�̷�̹���J�NFBMRAMKYJNJ[LA[GS[PO�N�D;C��_��       �[�&�F.���.pX(ٔ�ȫ    )(�����:X"(������W��`����7W)V��7 /W\�(7���@U��7����&��)�J�{���|  �����<�������t�'��G��0��Ϥ����0�����΁��o�����&����    �b�bF�b����)��J� �� �H/��"�Û�����)��)��K��)��&�&J>JJ������@�����)��)젰��q�� �� �?� ��@������@N �ȠJǨ/�Ȩ��A��o��I�  �
��Bȃb��b�j��O����������c�J
��

��J��0��d��0b�(/���(���(/������$� ������ӉlƁ<(�����  �����0 ��Z
���dƒ6��FȁL� � �

b!���
�9�w��A ����f�� �� � �(������  ������R��b��k � �l���������J����F.�໻7�J.
�����r��d��K�����&��B��{    ��� �  ���Á ��/�d���&�.�l�<!��& ?�/��֠�66
.

����������� 0֊KM?0C�4 �������4�� ��򈁂��� &!�ʀ����T)%D��E�X3S<ELJEF^%w·E�U����E��E��E�O6!&M66�BF�S6S\bkL�6����6E�&�FK�6��6GT7�'	F7]pA�ƪG�I�$ �NQ�� R��DL#� S`Q�	8�� �XUE�3 �  �D��ET`!�T@MN RP�	��0M�3����TN(�X�O3�8��D�X0D� �  OS� LQMN �P X�TL UٔCX��C	��QI�S�@1��TB	��QI�S�D1҃`N�@1SRN� ��ES�8�8GL��R�C2L	�� ��X0	���MBEB  � S� SB�TTNR`�E 0ٔCX��C	��T�ES� 0	E�O2�8�8G +�8Ne Ra��DN(MN!��CS� LR�1 S0��N	�8UE�3 T PS Um�T�RA�@TP 5Xm	E�3O�#`��B@ 0N%�L@̓	C�B@� 5�B3R� 0R��NB̓XAT�RL �RN X�@D ��3��ŔC R1T "�N �U��1��I�4N�!U�CS I�4T� DRNSQS  Փ@�P �S��MNQ 	S�H��C L�1 �3RT� 0S��?� ��ES�?8 R1T "�N �SO�X��C	���ES� 0SRN�`�BR1	��L�D`�� 1��S��`e����3� 0L#� N(�0T�@	�8�8G  N$ �Q8��C �Š#S�8UE�3 S(N�PO�#�մ��	�S�ES�	8�NEC� B@ 0O`eI�4LD�Y�� @L#� �R1N T҃	���CRT� 0N%�L@̓	C�B@� 5�B3R� PL#� ��TBP�`I	�c ��B@	8�S0��AD��@PT5D��3U�4`�N%Š�8A XS��	8�3�� F2	��� 5T �� 1R�MTR�U�4`�N%Š�8A OReT�`N  ��B@8S%����	�RN S�5��D��	�S�AC`�c8V`� FR�E�3�ET�HMN!��CD � �T@MN �Q�	5� 0� ��8L@!���"�����( ���"��k    ���"H����J��&�F.��&�F.��"��b� ���� ��� ��	6��C
�d	
7��J����[
�N0���