����  HA @ ��!    :  W<      ?  !             Z ^ b f <���������                                                                                                                                                                                                                                                                        �H�W�c�o�|ǝ!�+�G�Q�b�4�$C%��$�%")E8U8�T�cT�oT�KU�[U��T�jUxe<�eA�eF�eM�e��e֊e����h�U �]#GL*���ON(L`!�E3���8N`N$ �Q�4 E8L�s��&��R�t�BE8L�s��&O�tTD  ��3�Og�E�8T "TPM���XS�[D RL�s��&��R�t�BDRL���2�Og�T@D� ���E�u�QI��D`�8M@�N � 5ŔcRUuTXL@!��;U�TU���@8]��	8��6�4@rNR�(I ]G1LGT"	���d`q�E�8M�P��DCFCT O�# ��DG�M5N �B3RTX���n1 ���IsσG�҃�V�Cn! �M5N �Lg��2��kR���D��3��G R��C҃�Ѕ�HLn! L �0	�SL���2��kR���D L �0	�SL���2��TD���;I�8��4� 5XS. P�SN�`a�E��4�8��TS��  ]��8�	E�8��TT�`� ��2]��8�	E�8WE#L���2 ]��CW��	E�8L�	�`7���  ]��8�	E�8��TD RL�s�  ��;E�D��C�е��E��OB��< �N`!��R��T�5 � �T@D�M5N �B3R�    �A qR���A��4!Q � @      ��� �������������������
�T � ��'� �ŉl�(/ŖB��bF�����&�P.��/���� �� ���� ������/��)����ȟ��"����(/�𢯁���� ����� �F��  @G�� ��?@ ��`����_��`P���                                                                                                                                                                                                 ���v&xş                                                                         ��7�@ �� �� Z88��2�6����b_ � Y��� �B)�N��  �?����8���#�  
 �0  4���5� �8.����3���}��|��������?���+��04�c��~���c������/����6��{���l������z����"c���6��� ��z����,6�(?�Ѧ��� ��Ч�(?�ۦ��� ��ڧ�&� >�k y ����� �����������蟁��R#�P� �/�D�xÁ(���{)��x&�	&�&�Á	��J5�/�����l�<���w��b�|�5  	�&�&�nxb�bvi���u$�����/���i��� 	B�b�|�5  	��Á��tx���&��&�|�@�m��bf�ju@ee�@ BP�����@�o������4� �&�d���#f�&�)&sr��&6H/������� ��q %&� ��/�"#t��|�/�~�� �q �jq��s��(��p���z +���,(/�!�obun�u�Ǿ��si�p)��z�"�bF��&�s������m��j�&�b!�j�"&΁�'�b �j ����  �  B��~���� �&l9�k�ju� �� �� �� � % � > %b� %i �h&�&�h�(����bH����/�F�D�d��H��g�/�� �fbx&e&�ڈd(/�c�����J�J��K �^�+�Á���.b��b �ފ ���k%a"(��`�/�_�uv�^��0^k^�/��� q ���/�k��h��h��b�F��Ǳ� F�'�Ĭ��F��� p��]&x&�N$�h� �    2�o�u��(��!��mu)��Z��{ &!����� !\�(��[bcl�	&6l)��k�/���	�J���ȫt&(?���H�s �=m)<�&���;�y��/- � 0�/^#����Z*�\b�n/-f(?�H��|�����.����Y�!X⠣�+�/��q(�u�|0���W0t�J+�/�.�/O���2�j&!.obun�u��^�q0(��V�/�Y�u9U0TyCk�/��l����-�J-G�JS0���YR�u�S0����Y�Ru)y'��l9�T�ƒ� ��"��������������+b���X�+ !��n��4c(����/������k   ���Ĉt ����Ĉ� �!���c(���/�����6��� ���(���(/��(���@/��m"Qǚm&�o�Qn�Qě��$���ނ��d�����3���  @�����Z�j�#���� �� �� ����K�K�
Á�Ɣ.b��b ��� �����{(?������ `P�
�b�d���.2f��((cqO����(�((bN�/���(s0���(�B(+r���'�/�%�s��(� \�*f[&y0���*�N�J�*���@������� �!*�@����{����q  ?����~@�-@<�2��)�&(�&�!>m�/�ᢿ����&�!.)�/��!m⨋������&�!.)�/�(���cO�/����(�q0O�/���!.(�/�)��j��B!(����� ��(b(b�7���n&!.�/Ɓ��&m'(�D���( .\*&� �    �(/��kr����$t	c%� �)����ɥ��%� }�� ���<����í�b��f��0�����&��1�����D��� �᪠~��7��,�����&��D���       ��4�b�|�  ��� �����
&��'�b�f��?���j������/��ڠ���j��b�M)C���� �M)MM�~�� ����  �|����0 l�V��e������xÁ(��{��������z������������<zO���hÁ(υ�{)��h&�	&�&�Á	��J5�/���&�Á����w�&�,|�5  ƒ�b! ��k �L�    <aR��b��&�K"F�H���&�P.��/�󩀀�3�����G��&v��G+ ����4����>�b�nd�?����&�3�3'Ѐ�Ѐ�Ѐ�K�'��'m�'��'J&1�n�nIbc(���M)���
�"���1�&��� `����	�����3��i��� 	�� �����c�x@�`b�o��t ��܁�� � a	d����w����w�q�8�R;� �a��B�
��� ���� �����q�(����+�Á�ƥ�(�Á�Ʀ�(�` J
b`F(� � ��$�i�� 	]&�&� �Oͼ���k˼hb��b ��
ǁ�Ⱦ � �1(/�զ��� `��Pb
�i11b�u�����,��|��+|i�a�c�� �khPoH����oP�j ^��2�o���) �(��O�/��}�/��m����O"�j���M)� ��/���M���k ����M)�k4�/������������c(��M�������Ԧ�����*����Ԧ�����*���bM�M�����l &#6#\� .V �a�i��k �?`  _ g<�>���6 ���� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��D��D��D��D��D��D��D��D��D��D��D��D��D  ( (  �	
 n������ ? �<�>���������������� �%�&�'�(�)�,�.� .5	7[>{@]H}J^M~O\C|E_R � �� �� �� �� �� ñ �� �� ò �� �� ó �� �� ô �� �� �� �  ? ?	 ? 
  ? 	? ? 
                                                                                                                                                                                                                          �� �� �� �� �� �� �� �� ٠ �� �� �� �� �� ������)��)��)���n&�d�� �� �� �� ̠ �� �� �� �� ө �� �� �� �� ٠ �� Ԡ �� �� ٍ �� �� �� Ҡ �� �� �� �� �� �� ԍ �� l'	�} '� ���u��'�xR�k��� �  ��{�Ɗ��=6�h� ���Á�τ)� �� �&~')�J���s�@-�T���(�e�����7��D��J�����s���Ļrźy�R�pl"I�/���W��  %��U �%                                                                              