����  @       25?  ��������������������������������������������������������������������������������                                                                  �����2���8��ab�b�li�(/���)i�  �
�lI���cT@J
�cTJ
��d�42N(��6�+b�j��bc%c&c'c(jk(d܊�.	�li~r�vk�p� ^id�i�&*�,.�   ��(����n�n�liv��   ��lH�&P�'� ��&��� ��C�i� �;`.  � ���/�  v ���� ��� �
 ����g�����������������|`��   /0 :? @ �� � �                                 ��U��U��U��U �f�Vf.U$�f�� �u��U�J�� xIf ����/�%`�,D��E���&�^)�~����GfFDf��I�bI�/�,�I�/�;�IIb!H� ��DEb���3/5?&AOf?f"BBc(h�@iFD��@�D�/@o�(w�v(/�u��E���&>��O�J�����!�s��&sK�*!��"��*p'+o',�+ ���f�h���n �bD�.Hs�b �J��"�*���Ġ Q��E���'D�bc(��^[�#\)X��D�DD���BDbFF�DDbH��BDNDBc���π�B^9dݝBJ>JJ�7JJ
.k�Jk)4b)B
>k�Bk9d�_B�B�?�D�D��d�/��H�o� ���� ���7 �/^�d��_d�_�� ����� ���
�@.b/�F�u��#��r������ �e��LHbMLb�����bM����b)M�J_L��h�e3�r"bMrbbM��"�j"�M3brb)M�J"j)"M&�r"���8r"bM��_�r�J_h�el�B"bL�j!j)B70r�br�/�r���/�k�r
.k�rk)!j)B
>

�iB�Bi9B
>

�i"�MrbbM��B�L�J_��9r&���_h�i �Oy��m����U* �eH�MkiMO�3�bM��`��L�Lj)�b)`!�LL&�L�I�/�a�he��B&d�1H"M�bbM��`�RSfB!>LaiL�JBBC(��R%B@��S�nR5"bS�6b)`��d�/H"M�bbM��_�h�     e/�HM&kM����b��b;�H�/�)�M�bbM���)\)_H�M�bba�M�J`m�h�\3 2- OX e/�HM&kM����b��b)�\_�HM&4b)1b)�b)M�J_m�he��&"L&(?hJ�J
.

�KHbMJbiM���Ki)M�J`L��a��� & e	!L&�J&�M&��JJ&Jp)�b)M�J_L��!�L�bM�j�!�JJ&Jp)�b)M�J_L��h� �JX.XX�XK�KX.XX�K�+=�(�(�u� !��H���\2 e��L�bb_�L�Jhe�$L&0b)L�J<\) �he��J&HM&Jb)M�J_#�LHbMJbbM��`�L�JaJ�J+"���N N_d����PQfRSfNP$�@/���Q*B@���R$%@/�S��P�5b)4Q"b4�Rb)6S"b_�h��r��  ���?�+ ���Kr���� 	A�� �
��)��&�@���Ed�!�X�ec�b��e��JHbMMb���Jb)J-"�M�_�&?"���)\)�e�lB&c
�

�kJ�
�kJ�k"�jJ�(����/�J�bB70KKb:!.J�/�B�BBC���_��B
>

�iB�Bi9B
>

�i_��ԫ�����d��6� � z �ۢ�݂��d͊���  �������J� ��w)  J
�
��(��H�_��ee��B&�/�L�c�����LO�J�bJ�BJvB�JJ�b!B⨞��B��B&B"2���B"2���Bb9B�J#\)_a����<I"���ed�c�-�/�J�b_��=�d@�_h��*�L�nU �]L��g��*�LUiT�]L��g��*�LUiT�]L��g�������� ���&�yÉ
Θ���}�   �
����G�}� P��$�L�f�[iX��X]�L�Jg����]�� � �*L&YX�]�L�Jg��$L&[X��Y�X�]L��g��$�L�bCUi[X��Y� ��]��C[iX�� �]��LĻC�g��*L&�O�R��>( O�K ��L��g��]i� ��*�L�nOJ̠>�( �OS� ��L�Jg�]� ��ӛ�����ŀ�U�ԪĺD�*�L�n>( O�U�]L��g� �E�/�O�= /���>(/�O쀭�VQ̟��>�/n���[)X��Yn�� � �E�/�#��2b��n$�&1�&�H.��n�D.��b�=&>(/�=�!=� ���=�O��I��N�ʀ��󤷳�TܚW���J&J�'�\�O�/��� ��J���/qJ�� �     [� 	/��  �� ��� � ��� !�� �"�� $� �&�� ��< HJ���bƁ&��"��bƉ&��"��b7DF����"��bƔ&��"��bƚ&��� �   05bǛ �3b)��J� � 7 ��b3�8�"bԛ ,(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!� @   ���&��J��J��J� ���b��d������    ���� ��b)� ����b�� ���6��J_ǔ���

�
7�(����bȨ/�ȲiǓ7(�Ȧ��"����i)� � =?�"Ho���/o#�\_�ad�_�F�F��oh��R������Q�(�/�P������O�(�\���l)�� 0��f���
 9$� �=_i?�"!A⨀�N?b�A&dΝ?J.H0�k��?k)_A��di _	?(/�"�(��!(/���(���(/�$� ���Q�RSfIQ$*@/���R%B@��S�nQ(/�5�b4�Rb)6S"bd��_�aY��O�J�΀ �	�%1�>J�S\�lu�      �̼���!̀ �ȟ@���)�@�Di��o����Adp���_��D�/�F��@�G�/o�FF�ȡ�D�@�����FH�@D����D�/o?���/@?��?"���'?"���2�*�?"���D�/�3��(�?�/�D����5?&?f"BBc(��@@k �_��\Ҙ_ʛ �HM&�J&�L&Jb)JMD��L�J5J&%L&� ���V��U
	     u�����1���o��� �?�"���� ���F�F��E����T�����>( O�I��cY��O�J��=�n�?"���e!>��/�J���/�J��,�� ������b�mi��ǻJȹJ������� �   �������x���V��ʺ� ���i#�� �  U= \�p�)� �  D��!�k��� ��40��}�O ��#�\G�FOfF�F���F�F���7?(?"����_�ad����OciRRbbc�SSbbc�b_�ORb0FD?�S0 ??&?'"���?�"@���J���/�J������J� ��/�Ѫ�G�Ѡ�F?bfB&B(?�@�#\)@��� ��������� ������%��� ������1��� ����<���-�4��R�� �� ��������������������K ����� .��d��J��d� �    	�0  ��D  � � ��/�� �������'��; ���6��C�(�@��

�
���0(���@/��"ݔ� � RN�!�T1�C�. Ф� �������ïظ��ՠ@ �?p�/��   A �� �����;�������泲&�(?��������D�������)�)�������+��"��b8�&��6� �    5	>}�tq�on�m{�| �_�eF�JQ�k����g�ޛ�ݖ�y��{S��������d����� � � ��������� >��y�����������Š����x9�����	ef� d��������6�I��h� �   �)�9� ����������; ��/�����������TN"� ��m`���AN NB m[Ӆ�l�pȄ18`��.8G�נK m�`�ŠT�D8S.   ����8�� ?��"�����'��J������ ��.��pݧ�W> nb��df�e/�� 	 �� �����/�����)�)�Y����b�i��F��6��J� �!�⨶���2Ȳ���2�����0��{�)����� � �
   鐨����6쐠��#Q&���P�n$N&Pm)�r�N�JQO〮�P"PPb�H/���m�〮r)� � 5  ?� Q��PS��HP���/�	 �N ��`O   F��b��b����d���    ��)� .��b�����  ��y��� ��|���|�������� ����7r�8r�9r�:r�;r�<r�=r�>r�?r�@r�Ar�Br�Cr�Dr�Er�Fr�Gr�Hr�Ir�Jr�{�����w��f��f��f��e��Y efd�������� � 	�I����c� � ���/���&!̑"������ �헲����    ���������b���������P�X��Z��]��`��ȟ����Ƞ���'��	� �LD �N�� z @:� ����� ������ ���&��'�H��ϑ�������� /�3�B�FCDENF�	(�X��H�	HLC����2֙CW�؁Yڕ@[����H_X?��
8��H � J&!��%�� ��� "V�"��" 	3  �  ��3��3� 41 H  �  �  �  � F�PZD��D��D  �  �  �  � Ʉ� ET� %�?K N%�`�R C�E��O��3NB�P`�RC �T�T���AB�TR�5�?K UP28N`!�DS�? PɇC8N`!�DS�,�_�� �C@`�?K �RN %�T? �NB	�S��UNA��PQS�? P��@�8E �T��N%��@8S? 	�S,���RC �TCS�  PL NB�P`���3NB�P@�RC �TP�D��2B�c� H�S`�CD�4N%� @	�3Ȁ�5� KS� �T P�C��8�$�R�	�8���T ��5�E ��0�����@R��R C��@���T ��0�����@R��@BN2TO�8(�@1N NM1�C2L� �0���D1����0DT�H���T ��01��<���RC �T���NBT`ԉD�8T "`� C[���NBT`�5TXT "�C��N$ �S��T��C���DT �4�N�!�LC	�S N��2��@C[� ��Ȁ�5� @�	S �	8��D�Q S" ����M5��; �N �8S��LC �S 8NB�P`�RC �T����0S� �SBR1  �? �N �8S�? ��TM��� ��  ��N�4 S(RI� 3SNR�O-�T �� �T�4��E �	G��4C(L #�N?X �	��E�NBL�6 1���O0��CS� U�NBTD��H�8��CB���@R�8S%��1��@ 8���������� �� 5N���M5�8�8S ��������/�������������k   �L@8� � HP���	 �
� ��7ݡ@� fhg���� H����Y0��s
����"��y�A0��~��y�A0��&q .��b����Ӛ�E0pqbD�!p⨮�p>"4p&�?2 �c�op�  r� &pE ��bH
���& �0� 'p�&�X� ��� &p� �r>�&��J��Ā �� �s�� b� �q .if`g&�㸏E X
l ����n�op ��@��U  �