����   � �   ��� @�10(<H 2'?!	  ".2'?'  ,".
-2,,22'?!! 8".>2'=2"4242'?"   4".2'?*  9".2/<!   >
.;...I;?::<$ >4>A;''2 ??�B B <���������                                                                                                                                                                                                                                                                      �� W                                    �!1@                  .墼��                  �5 �                                  �	Ł��� � ��<����b�c(��	c(���	Ǒ�ʃ��*�<�� � Z	���  � � � � *��(ϫ �Z&�!�� > �   �j/�P�t
                        s��O/            ~�.�                               S���(� �8  ���&��i�(���������(���(/�@������i�����(/�������|�@��"��������"��&�*��b��������&��/�����d�����/˃�~����n��b����j�H/��� �����/���}��i��� ���|˃�˃{�          8 ���Å�q����� ������K �F��� �                                                                     �q�                  �%  M                              Ӽ� P                              [qp<���I ������ �,���,��7����A�K8������Ɂ�ȁ4ǂ�ɀ �4���Ɉ �9����P�� ���"��k            �1�                        ��#*#      ؗ J�                        � �                �� 鴇�                        �!V@            �  �                                                                                    ���      �e���                                                                                                                                                                                                                                          z��s                  e�0�G/                                                      N   �                                                 ��  �
      �� 4            es0 �                   8  j� �� 0                   �	�Ф�����É� ����'��&��&��r��r��y�������k|����� ���n��� ���� �� /�/��!��&��)����L�<��{ �	���׀��������ـ��Ls� �ң? �P�	�S����5 �A q�TB�  P�	�SB�GO%S P���� ϻ�T����Հ�P��Հ�P��Հ�P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P � L� �&Q�#A������#A���PF0�#A���� 4�#A���	 S�#A��� 0�#A�����#A�� 0�#A�U�T  �#A���� @�#A�E�@A�#A����@�#A��DR�#A��T�#A���4�#A���P�CD��8 0�#A���F �#A��PP�#A���TLR֟I����#A�����#A����#A����#A����T�#A����T�#A���T��#A��T�#A� �Z _��T����Հ�P��Հ�P��Հ�P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P��P�c	.��Jq�E�k���j���JR�`��g	k.wׅ4z�ޯ�|h�l���צ��[n��p�A>��m�D
֒��)��A8Y��,P������� �8��@s�t�ۗ��!t�Ɇ^����Q�V�ӿ���-����?�Ѭ��h�)�)�2���� :�8�=Q8����nlyS�b�ԃ[��ư��                                                                                                                                                                                                /,dD	�J�VT]�է�<�Ñ�p��H��k�
o&��K�Q���N�O��tf�Y?�s��k��"�c�$��X���s�q�)����"`mYg�cM��A���{��ZRԖ	::[������̼��Ah�FL��@��2���<q(\ߌ�+�pڲ_�������5FR�啯�D����R$�ߛ�fv�n��a*�٥� ��DW��G��dȾ��8�oIO`GK��%h�!�����r��c�y�����kN P������V"E���7��Q^T�?��<6���	�ߴF]mD��¨}�ދr�(��}3�~n��ֹ��w��8�VҖ��!��^7�.x3a>u*�+~۫J_~̊�?K/LO�డj�أ9�:*�f&Zǆ�������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc�������(|R�¨�����D�뢠����Ɉ ����D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ����'p�  � 8 ��}���v	P�nݏ_��Fm n�&8H.�����H/C�/�ڮ�/����"�i���&�!.��/�Ȩ����}Ɉ ��b�bW�ԉl�@�|"����"��l�'����"����J��B(���}Ɉ � ���k�HB�?�D����Ի��g?�"���V�"�����'�N��PTB 0��� ����� � �,�` VV�!�۠/�F����۶��r��x|&���(��m�/����(��m�(��@��|&��y�����m(/��������z�� �"�b��F.��+�(/���H��bV���������m� ����⨉���۠/���V���(����������`����? 8����W�f'2��pD�F�&�`>E��� E��
���	&u&A�.��&��r��/ @��f�����|�&�J��|�&O������ݨ*���C 	�u�C !��H��	�r�A��F�?����r��	�'|�� /����"��s��{����(?��B6� � �� �  ���pWgJ��(���o p�x�݈����/���}�� %����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ����� �  @���     8bD8��&m F���@/�ԦP���J�כ����O���������� �v �  ��� ��0 ��� ��(� �&!̑���������c���J�޴�����2X��(?�
�

��������ς����o��R1��D��� N E��D� �@C劀���	��T P�ل�MA	O���� 0���/a�  �f�	&�	��J�g�v��KV�e�� �@� �? ����   P H  H H� � @�10(<H 2'?!	  ".2'?'  ,".
-2,,22'?!! 8".>2'=2"4242'?"   4".2'?*  9".2/<!   >
.;...I;?::<$ >4>A;''2 ??�B B <���������                                                                                                                                                                                                                Q8V��/�8�������m�(��@��|&8&8J.8����(���H/�J�V�8&��,� ���S��'�J>
��H.��J
��������u��(��!�瘨Ϩ �  � ���J^
�?H.��J
��� ��J.8��8�c8V�k              � g�P�@ ��� ��\�_"VU�2d� p �     �       �       �       �       �       �       �       �       �       �       �       �       �       �       �     띓��@��������Ӎ� ������?�!�}] c��   ��U�����D �B � ��                                                                                                                                   	 	                                                                                                                                                                                                                           � ��G��"����Z� �	�����  �	�Ԁ��	�� �� �� ��  (����/�ؾ���(����������  �   ��6��C�b�����2������    ��F���b���k �	�?����{�O�MN0 �3� 0��[               �T^���?�
G~T�����Z  ��������� ���|����� ������7��������&��2����Κ� ��㚣 ��U�� ��ۚ�ӳ�-�����-��� � S	Ut�DAN�!�R���DN(�A3� 0BT��QIu�NB�S�n �LS!ЃE:! �LS!L�TD� �                   �y�c�VG�V��?�������FN���&��,��|��C����������i�����i��������(������I �&���� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d��������D��� ���޴ � (����B���ǉ������˛���������� 5�����(���ɀ �5���K���< ����F��C�A�s �TEB3R �ϋR���DIV�8��4� �A q��@C1	�S                                                         �(�Ӏ��? ��)��7�����'��'��+ ���bg��J� ��]�R1��� 0���R���D�E���PL� �?�4R���D                                                                                                   ��:-^���������� � ���� �ᆢ��b�b��ǉ�Ȁ���<(����b��/��������"�������&�����* ������� ���ǉ����/��� ����  ����ӇD���&���ֈ������� ��� ���d�(?ֲ���J �	����$��+ �            � �����`�� xE���/�������2�����̨�� 7�����2(����/�����~��x����� ���ɀ ��� �� ���É����������'��'����:��̀`Sr�݀��0�H��A�3�N�G`����d� Љ��Y��A qO�3�T                            ��������%�V]y������,������ ���Ǹ��b�ψ������������� ���F.������&����&� .��&��"�Ղ�&��)���ւ�������փ����D���� ���&��(��J� ��р�� �       ���"��b�ڋ                � �@�?P	������S �U���	B  ���)��)����֞�����)�����)�����������	�����O~�Z<�? BYPG�                                                                                                                                       �  ��������� ���Ɂ�́����,���������#��ǂ�ɀ � �	��ɀ �6�	��Ɉ ��	���  ��	��Ɉ ��	��ˁ�É���ǲ��Ɂ ω��􃜁 ���ɀ �)�	���	 �0�	��Ɉ  4�	��������< ���� 4 ����� �   O��?�u �u8�� �G������&��&��tφJ����
�C � ��'��^��ǉ��8  ���� > ǂ��H� N ǜ� ���w��|���� �>����H �N�σ������Ɂ ΁��� ������&� �   ���(����s�����0�/��͉l����H�����@ u���� t
xG:� ��E��������������                                                                                                                                                                                                �   �xş          �              �                   �p����d�ާ�و���������8����� �k�Z��O� 	��?�?PPS�������_K�λ��t*�F�	��	 �gP`v� v�s@�
܁�*� ��Ƈ`�D� Q�;�U���u������!>~�/�}�����������|y{z)yxrw��v�(��ui�9�{���ô��� �'��q��� ���ⲇ�{ࡨ��G��4�1�����,��7�����k�� t ��4��c� �qc��͒��͛ ��pb�l�.����&��� ����'8� ����/����tہ������ �0i͐��7g� ���g�&o�ui'�v>�s7�eI�I�I��q�}��kL� Ө/�n�'��m�/�l��zY���&z9��|�wk&��Kkr|i{z)(?�z��{�z��jz)i"z|�� ��f���Bf�e�F�&h(��d�(���@.c/����b���� ��; �&�����퀕 b	a`��r� !�/�r�!�/�΢���r �!⠂�r�!⠂���/�r����� ���b��f΀h� � ���&��&΀h�|�_D� 1^{ ���&��&���ċ ]	_��8Մ3 ^_Ο��4� 0^{_��L !� V^�����     � p� p ? ?`��؇��    \��b�vi�/�����?��[�/���b��i�Z�     ���v���)�/��b(���b�Z�  �
�Z�	�Y�y���X侓��W�@W���/V��bU�&T)b��rc�&��JS�"��b!�����@>Z�/W�!��!.�?W� ����J��w ��p�dtZ^3Uf3u�����/R��^���/^R�����r�؈�_ӟS `^ ���'QP��u�C��T��F�� �� Q	Or� !�/Nr�!�/N��uS��T/�C/�  �M�R��e�r�U(`��/��L�r��s��_��� ^[ b�kK !��hK��/�g��J h	�j_ğVC@^y� 3X� r	Xs�� ��QiJ��r�Is	u	S�T� �K !��hK���/�g�A�h��j ��(��HZ�kv����(/�[��R�&&Q�b b�R�^�^J�r �riå���r��{�Z�	N �G��Z���JyF�pE)�ρ �r��riH ��+ 6/"�"H. r	L	��J��"�e���s�s)^���QP����MR�r���@.�/e���&Π/������D�zG�w��M���,�^{ �q�"��b�QiJu�C�� Ѓ RM^�s)^r��D�zG�wК�ۨ^ ���Á��� ��Cb��b�U�z����d��   v����_ΟM@^0���"�b��a`��F�!!b!"⨔�|!�"�h�z)r����z)ք� r	 �	r����z���r���||�_��  �)�)�z)�) �)#(/^T���&|_�υ` �^b�a`��r���r�Ȝ��Ȋ r	�	r����z֛]_��^� �։lց<$��� �SE)��ā���B)g퀸� ���	
�)_ȟNR�^ ���s�$��c��{   �(?���������J��Ck��������� ���6��C��d� �   ���_ٔ�RA�O��� Abg�J� ���bH/�!�w�/ۼ�"��bZ�����,�_�ω�ɀ� �ZB)  ��B) 6 %�/E)� ˉ ��_����@^���%���ؑ�gvQP�uF�	 X PR��QO��&c"�b�F��ri�ZZ"�b�&!.�E)� �� ��!.&�&����bT!��bc�&aʚ�F�a������r��s)�
c"ܶj!.ܠ/��!��&`ך��!��E�� � �!��&@y� ��&� �(/^�����R�����?�����2�ET��� ��bfJi�_��� P^ �~'?>'�='Z�'��~��~<%6��������j��JK T�Ӡ��bKt� �   ��鵠���b��b�d�Ӫ��� ��;³ff�n��n��bhi(��b�@.��/���@.�/�u�R�� �_ӟNe ^k_ğ� @^��P?� ���E�����D�&�&����b	�b
�b�b�n"bia`��r�������� �F!�!""����rI���!!."�k��r�������!'�	�r�rib���.X�
'r����r�H 'r����r�J�s������ �q:0J�(���ְ��fـfɔbF�t�����Ѽ��� �"����+��^��y(/��&& &Or���r�Zs�� r	T	U(q�F�ri9 �+ �	�!���x��������'r����r�H �'�!���w���?���8r��{�(� �(��7L)ri���r����V�j�������������� f�U�u
��_ZB) �6?2�5c?�&wB) �4E)��ʁ�4E)��ʁ�EB) �3Ų����B)o�#D.'�q�rU�&2E)�ρ��E)��ρ���Z���&E)�ω��������$�c�9���i�/9�"��x&!.��+ ���'�F���i&�ir���s��������pE)�ω ���7��Z���8ZsjY���m� ���l�����6�,� � ���Á�Z&�&@y���Z	�� ������7��7��r��ǁ��#$���!.��wn�b �� �� /� /(��C�(���(/��(����R�)b�����J����#6�#+��B��z��(�2����"d!)b�\�[�&������@�� ��#�qG�/Q*@r��92;o c&��@Z☀��C��� �!>��i@>Z�/����� ����c���b���?��B �?	1�( ���1�(��)�1�(7����?��B �?	� ��&��6��&X�B �?�B) ?Ǜ r	T	U(!�ri(/���!�:�&���8   �   _��� @^���7a��4�E�����p4E�����'�	a����.�cE���� 0�E�� �� ��b�b	c(���	cT/�(��µ&1B)��J�	�� ��à���M�9�e�� �����/R�#^k��/E)� �� �3B)  �1B) 6  .�E��'��$��ǁ_���D�L Y����@ ;��z���T ����c��d��6��C��d��6��B����������D���� ��,��/��� � ���9��<�p�qK��?�_��TR`��HRC!? P9w)�v�G ��/���� �F��� J

�� ���b����&,!�ʀ��� �@>��/��� � q'�彠����E�S����Y� �E�x}� ��nc���J�?�������� ���)������ � (����b�¨�����"�����Ĩ/��� ���8��4����� ��)��)ށ���{ �	!��܁<������D	�T5 ���Á��� �s  ��h��)� ���$����)� ���f܊ � (i��� �q�? PU��  ���样⨟���&��"��b��l��6��É��ё,��t ��􏁬��&��"��b��l��6��É��с,��t��D�����       �	��D�����  ��Ǥ��&��&��&�Ѫ�ߪ��&�0J
�
.
���󣚹��C���ȯ�������� �� �      �����矣����                                                                                                    �-�<,�/�+��_�D0�: ��ˊ����|�_�D: ��h׋�������^ �*w)������������w����*�� "uˮ ��X�q � �C@S �� � #��@�P#��@�$ � υ � EO3� @˅�OB � �R@ �P��%�@͌ ��2�DN � �$�� F ��F �� � ��0� 0�	� 0�� @͏	�4 � �T2 � �A3�  υ� E�A@��OC� P҅� � �� @ڏ� � X� 0��� �UP2 � �RE �@MG @�U3P  ��R T�� � N�%� @��F %�� F � �P�	3� 0ŏ� � � Ǐ�G0 � ��0� 0�D  ̏	�4 � ��3G  Ϗ�TC � ��4E 0�� ���LR � X� 0Œ E�!Ɓ� @�� � ��0� 0�� ��DÏ�T0 � D� @�UE %�� @��NB � @V�NT � ��TO  �2���	�4 � �# � ��C � � ��R Ǐ �  P�� 	SA � ண � I�	^ � �$��� L '   � �� `� TR��� Z�	^���� ^�� �  	� ������£�   q �	 �� `��� �� b�� /	 � �|���� �����ض��  ���9�� ����?�� ����<趤�  b���� ്� ���ʎ �� N 

�� ྍ�	 � �ί�� �Ϸ�趣��@  b��� �г�* �� `   ! � ��� � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                