����   !'==.<(.!'=*"M= N   ,?".   
89: 	?=	0
".    >"=".  0&0!*; .  <7;82"':	   
78
8" 
8'9".    O9!  
0A, > ?  ? < ? 8?  > >                                                                                                                                                                                                ϖ��@v&xş��C ���G �                        �&���(ˁp�   ���8 �t�C ���0���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�?� @� ��8������������ ���������։L~/}A?P
�
�|6{6z6y6x(?�&}�<������lw�<������lw�<��  �	�&� ��$���*#�/��K y��  
�ظ� �x��  `���O �� ?�!��� 
.

������ z (��~z ~)���R?�y	� 
� ���� N�i� ���ܓ�bv�&�����4��cuD!���4t��!.�/�ޢ�ޒ�b��������������)��2�������&�wÁ����  ����	��ՓTUL�`� 8�)���0� @�w�  � �bi ��Xp@��u@ee�@ B�S!3�1 � ��!��"�� �2 ���J$�i� 	 �
����b��c��Kh����� ����i� T?�
����  �������̀@ �����d��2����ӊ����P.��/�٨�!���0��O�٨����J�ъ���ǀ������?  ���J�
>

�堮��c��@��b���� /��@� � ? ?`��؇�� �  � ���b��k��b��k�b��bs.r�A����Bs.r�A����D���F��  ��w���b�d��� �                                 �2@G�"o����""�j T F��{'�+��D. b ��p�Yb!�l!tF��!�zE�i� * 2
" ����q���d���(��� �p�Ao��� o��� ��.nb&�)�bn"b��� � �A��)�@��?)u��>&����B�/����)�) &�)�����4(���/�פ�ף  ku�D)t&(?���H�s �=m)<�&���;�y�� 7 � ��S��oB�R1��DT ��(�m� .
�����
.���)� ���4�A�n�(���A�n(����*��*� pਰ�v&xϐ�	HA�1�� 7|>�������	w�k�x�ԃՃ� 0 �8�8�8����D7)8)���|ly���a�S��*���{�x9��E����3 l ��(� ���bD��Pp�(� � ������� &!����� ���c��l����R@	�S���D ��
����� � ����,�'��;�� �i ]��J��'! �����6��C��b�(�o������ �
��$���ނ��d�����3���   ����   J
�
�!8���� 