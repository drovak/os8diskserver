����   � �    	 	-08-	-     |)B =+��������������������������������������������������������������������������������                                                                                                                                                                                                                                            �8�  ���L !�Lߌ���fE ��ʛ5                                       �  �8 a   @=a   � a	            ��� TP P�A[�� @ a �  J V �A R @��A �R�  P` e�             � �A �@?� �	�������������Iҳ���É�Ɂ�É��Ҡ������������ ����� .��d��J��d�\�   � � 	��@ � H �� ���É�ό��ȁ���<� �������'��; ���6��C�(�@��

�
����0(���@/��"��� � � @�?J�H�  ,�!" i ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}on�m{�|q� @DLZ�]��g�ٛ�ؖ��y�|ˀ�ؠ/����&��I������   ���������   ���q���� ���
���kƂ ����@�JIH"bc"ia"��������6��H��h� �   ��)��9��� ��?�>��� �������d���������� �	���/������,�<�����Ҙ��<�|��&�Ҙ��ÉF����ǉ���� !�/�����/�����/���������k   ��H �P���>�I   H��iac"b"HJ"� ��(����@O��i��� �F��b��b��ʜ�d���    ���(� .��bʫ����   ���A������������ ����� �	�ɔ����ɆȾ+    �ߠ/�ޢ&!��"��ޢ��� ��ײ����   �������TRN�!   ����<�����  �Ɋ �� ���� �	 �� ����� ����� ����� ��������������)�����)�Ē��)���ȱ�����ȟ�����y����	��C@ ��LD!  ��N C�� �Q�> �����TN"������ ��׊ ����c��{ ���É����K �	 ��� ����� ��� �����?� 2�1����� ��� �  p   ��!       �L ��   ����&��"L  d�����RUY^c�����TV � UB�v� C�]$OD���e��i��̀�� @    ���� �������
 <����� �P�   ���                �� �   ����M�                 � ����y�i.���?)��wyDfuNbI^fd�nH�nG�iB&�%�������CJf@>��.���(����wD�n�NrI-i\o&P )����o�������o2i�a��)*��4���?�}�!�����3y3��=����g�"�����2���� ��@���V �k��|�*[�� ���D� L܅� �I��Z1�K3	s��.�ei�����}b������"����/���b!�����/���b��/�������!.�/����e J
�
����ne�Hz���6ə���������R��U����Y������K^��޴�c������Kh��6�2������ �S�F J1�I�L����L�/��&W�*�/�/W�&��&0-�,��A5�p�J9���0�-���dr`�k�A�6p��*��0�-,��6�p�J9�����e� (����/�Ѿd�z�kN�Ii����ct��I������+re aE  3ޜ3*���� 3	g�ܔ�� �@�� ����+��@� �P !����0@��8U�A65���3�����#��c��k��!�"eF���b�vf��z���"		b
�b��r��{&
"!	� ��d�*H��_��	� �v�a�|�j���v�|�j�|�v|"v	d �������"��"ր.3�<�U�V�)�;�ee���z���&3e�� �@g���2���牼!t��d0��U�Z��o� .��f qA��.[/i+���&\n&\o&� �����$��|�#��oO����o�2͞\o&�z��!�n�������n�jd`&_^&�D>��)2˞�]����n�/����/��&�����3� 	�.��2��\�n�cD���j�������ijf���i�����"��{�� h1R3�ą�|ZS 뜺&B�* �>[/i\i&+\�jmfklf\n&\o&��!���aࠣ�nO����n�2˞�[�����F�(����mI�����3�Ḻ3�3�ȟ.��m["����F�(����d`&_^&�D>��)2˞�ߚ\!.j(/�\����2���[����l�/�j�l2i���m�/�j�m2i���2Þ]�J�@�9 i��h��3����a��\bo�i�� ���F���i$��'"�b��&��zJ|/U!�/��(l��k��[�/�F����l�/����3�Ẻ3��/�3��º3�3���&�z�����&3��3 �������F����3��
!.	&;�:���zJ|/Uw;w�:
�;�F�K      �+�h��t&
$B3��=�3\����'��oO����o����z�J��U��y��F������?���3���?�3���;�F����3�;F��2��F�(����ȟ.��D*I�Ĵ�G�Z�/��"�Zf��)�����3��.��ě�]�y�/����s��d�y������6yl�o�����gd $  )�@�@���s��3��B{�f�(/��&�Pn�.��b���(�(O���� .���F.�怽���"������3D�3ޜ��C�/�3�U.�3N�C(I� �  �    �� .����"���3"�;��3,���/���4��]�np�b����ٴ38���/�3�&ٻ3B�-;��*I�٫ ��NbI.i��t�JI�J��+��K��f���;� �S�F��6����ZB �ppb!q��d`&�e H
���&��&�*�*8UA�U�eU�Q��'��'���d�c��c��j��!qp"����*d.�q�p�/���d�Kd&!.d�/�d�!����:�=	���ՅsCa Q�1L	�� qp�/큮p�p�Np����qp"H�뗑UV���f�b8�qp"���pA.p�p!.q�jd!.�/�q�pH.!��d�kqp"���pD.�p&p!.qb!�p�/���qp"����p�p!.qdb!��(�d�k�_y7i��S��F��6�K���n��b@H����J��bY(��W�&��"<����JT�J��/��T�f��&���<� � � ? ��j�ఠ8AUJ b �]�f���f�[(/f�Of�Nzਖ�ffD� /f.��b�H/�����⸸&���_b!_����_!.�/�d�D�_�r�k k���jk&2Ş�N���@��T�` I3T�;e�3�������"��������"���3ϛ;�3ӛ;�3כ;�3ܛ;�� ���,��s���HL.���j�����7i��f��‖6��"!��h��!���B<����� �@Қy�/�����F��8��4��� ���` ��y�k�(/���@�<������j��hźK��(��(��&����f@Қ&,�y���yO�L�"��"����۶����F.��b
����bۜ�� @i����X� y︊���@;��j��H �n�l~�!��y�/�"��D����D�G�Ͷu����'"�Ua��2���QE  J����z�a �� ��%���a�������)3לD�bD�� �   B�s�H.��&�(?�!�\(/숯Q�#��6��Z1 �K�Z�b����d"��&��Z1 �Ko�����K��MM�i?6�w�; ��w@L��r��v �D�i� �D�J�D�D�k��̠���s�����2��e�1� K ��2%i ��Ers�b��/ꅢ��/�Q�B�&%� "�Ub�P2B�&%� "�Uc��a ������� ���b��J��2��e�1� K bH.
 ���b��J��2��e�1� K �����
�E[�K�K   h h]���MBŌ�~�@[ �� ?H����3��������F�/�����/�3��3���������/�3�ʤ����;s�:���2���;a�:���2����3��:�3	�:�3	���;b�:�;c�:��͚�֚^�/�3��ֺ;`�:�;^�:!�����2�����2�����2���3ƛ�;�d:	&;	_:	+G��� WVe�i��MB��g��g�����b�"(��N(/�M��(�ȟ.c�������E�E�-����E�����t��N'�����E6��z���+���E)��'W�&�'�$��_#)$��d#)�Һ ��a���oO����o�2͞��&�!.��2�db!`���^�/�d�D���d�D���          ����ʾ�@���w��@� � ����[��⋋e�1�   ��uub�ލ��B�&%����^�k3��3�6�è��3?���"���J3IDZ¨��3M�}�'�4y��?���3��;��3�e3�j;�C3	m3ɉ;�J3	s�˜O�7O���4<��G�b���3 �Hi���8�������� ��y�� �W�'�ٵ��;�x�@pj�II�d�|O �W3���
&-���&3"���2�8i�3	��(?��;�:�Y
"ȡ�3A�Y�Y
"��&��&3 �3��
�J�D>��&��"�3i�=��3ɚ=��*ɂ����̣���̱����?��K Ҩ��K  �� b�����X�Qn���b��@  ��6�>��nT;i  ���K�� ���°���O3|��&	&��&(?�?�3�����w&;w�:�	w6	x6=w��	"b
c(��:�
w6
x6=w���"�&-������"

bc���:�;��3��
6;�3��*��	&��	�d�3����Vy����@֛��������dg�h�L�&g@.HP����g�hD.g�+� ��N��M�M ���D�FNI&��2���3\���.���(����&�ߘ���� �b		c(��bt�����s��sMw;w����k�S�Z_d �y�/���3��;Ú� ������ /�y�����y��ﲠ���y��׺��2�����2���3͛���W���s�r�
��eg����oq`��G;wV�����i�� @	����K��&�̺�ɀ@���� �� �����6y�/��� � 쐀N���� �Σi �Mq�`1	G��4C(S�"@Qĉt��T�C�D� �  ��qVS!ԃ킕 L� �4�R@ XL ##� p�8vV�C`!�	�� �LC 	Q�TAX��E��GLC U�HRM TR��G��4��AS T ��� p Ň�8�� H	�� �D ���7VC`�HN�QT�  ��p�8 ă`�`@�� H �R�  XS� T� @��c] NT" �@�g�=8 	� ` R�$= �S� `_ ��E@ҷA- ���T� � �N  T` R�� @τT �  Pσ � ���  �ST�`R��D�MuC��	� @� 0��sLD= ���	q�TAX��E� ���DA��`5� @��tTS	�P 3���T�5(U�AS	�PP@�S�B� Q�u�HRM TR� Hߕt�	5E=8 �S��D  � T�STC@	��R1MXP� P�uC�C� � HL��  R���D ������T���D�` �/ �@ҵT@!�D@  P�8�HTXT@ �KA �E ��C� @�SrɇC �A�4 ��6C R���'S�$�8��C���N�Rנ3R@$�Ip�C1p-�	��    �R1�� �DM�P��HG1L*�����D