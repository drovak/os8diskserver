����   $<$6  : /?  0: 
68
799*+8*)2>222:'=.$?9        : 2>8 
:22:/<  : ? /?+<>9>//;g;55 29'������������������������������������������������������������                                                                                                                                                                                                 
 ���� ��� ���L �   ����� ������� ���?      �U�]$8�ǪIm+���ސ:Ԋp >���� t�W��? �� ?V�R��(V��HZ� r�K���Z֩A�?����s�
��� �v���? ���?��~z {| }���� *� o� *!�� ��+� o+�!�� ��� o��  ����& �� /��,�& �,!.� /��-�& �-!.� /��.�& �.!.� /��/�& �/!.� /��0 & �0!.  /��1 & �1!.  /��2 & �2!.  /��3 & �3!.  /�� ����,  �"�!� ��� "! /�� &_  /��z!>~ /��z!!~� ��z� e� !.z . ��{�!z� ���{!z /��{ &_ �!{�  ���|!>{ /��|!!{� ��|� e� !.| . ��}�!|� ���}!| /��} &_ �!}�  ���������~�!}� ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���e � . ���a"  � �  ��a" �  ��	&		 . ���		a	"  ���	&		r) . ���		c�	�' . ���		a	&"  ���	&		% . ���		a	$"  ���	&		# . ���		a	""  ���	&		! . ���		a	 "  ���	&	 ^	"  �����!����H/��		a	"  ���	&		 . ���

a
"  ���
&

 . ���

g
)"  ���
&
�>
'"  ���
&

& . ���

a
%"  ���
&

$ . ���

a
#"  ���
&

" . ���

a
!"  ���
&

  . ���

e 
� . ���

a
"  ���
&

 . ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���e � . ���a"  ���& . ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���e � . ���a" �  ��& . ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���������3��e � . ���a"  ���& . ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���e � . ���a"  ���& . ���a"  ���& . ���g)"  ���&�>'"  ���&& . ���a%"  ���&$ . ���a#"  ���&" . ���a!"  ���&  . ���e � . ���a"  ���& . ������&�����/�!^� /���Ri��/�!^� /������	� !����& ���� _ �!��� !����&���� ^ � !.ݠ/ �!π��b���� ^ � !.�/�� o��� !����&,o	f � . � b!��� !����&&�"�% o�  �� !.��/ �!π��blO<�? o� � b!��� !����&��Q�U o �!��� !����&�d�g o�!�� � !.5�/��� n ���T.T . � !����&,�f � !.��/ �!π��l!���� o �!��� !����&�������������!����"���& �  � ��o� !����&����f � !.�/ �!π��l������ o �!�����l �  ̋�	|���0 . ���!� ��?�� ���a � ���?�. ���>�. ���0. � ��0� � ���?�.0 . ���0Q. � ��0�Q � ���?�.0 . ���?�.0 . ���1. � ���1 � ���?�.���?�. ������ �� ?����~�{��C �������{"� ?����~�}�� ���瀦��� � ?����~�X�H� ��H怸�T( � ?��(�n�P�� ��� ��<� ?�� �n�8�& ?���n�/����������k��.��b��/����&,!��� �	���1 . ������� p��@�   �&f��K �                     ��"   LG�2                                  ��"� P�D ���2 @����ͻ                                                                        ���	���� � �!��!��� ���� !����� !����&� � �������&�� ����� ��4� ����4D �� �4� ���l4� �B
� ��������l� � ��� �� ����n� ������Y�!� ���� ���� ���� � ����7� � ���� ����� ��)�3-� � ��3�/ . ����� ���� ��`���`��<�`(����� ���� ���<�/ ��>� ���?�/ ���P ���P��.�P��.‡⠢� ���/���c!�⨗�!.��/���� �&�'����6 ���� ��⸷b��d��������&������� �    ����� n��,��� ��/�����/�H������ ��.��� ��<�� ��������</��</��<�/ ���.�/ ����P@݁��