����   � @         - 	       =  : - 		        01 	  		    	 	    �&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{ �(?��B6� � �gWq���� g�t��D�8�  ���L !�Lߌ���fE ��ʛ5                                       �  �8 a   @=a   � a	            ��� TP P�A[�� @ a �  J V �A R @��A �R�  P` e�             � �A �@?� �	�������������Iϰ���)��É��Ϟ������������ ����� .��d��J��d�n�      	�m� �D  ���� ����<Ȍ��Ū��É�� ������s� ������d��0(��@�
�

����(��@����)��J       � @�?F�D�  (�!" � ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    18}on�m{�| �>CLTb���y������/�������v��y�|Ӏ��/����&��I򀘀��   ���q���� ���
���k�����Z@�FED"��"��"��������6��H��h� �   ��)��9��� ��?�>��� �������ǒ������� ����岠����I����É����)��Y�����ǉ����iс��<F���<�|��J� �!������2�����2�����0��{�喩 �   ��H �P���:�E   P�����"�"DF"� ��(����`O   F��b��b��Ƙ�d���    ���(� .��bƧ����   ���A����������� ��� �	�Ŕ��ņĺ+    �ڠ/�٢&!��"��٢��ر�ڲ��� �   � ����J� �混t��0J���&��w��D�� �����"̊ �� ��� �l�Ao��n��&� �����?�����������)�����)�����)�Ē��)���ȱ�����ȟ�����y����	��C@ ��LD!  ��N C�� �Q�> �����TN"������ ��׊ ����c��{ ���É����K �	 ��� ����� ��� �����?� 2�1������  �	����������	  �5������ �R  ��� �E 0��� 	@3��� �BR1 ��� U`A� ���� @��� �Q8VC@�� υ	A�� ��� �QN Q�ȀI�R���H�8T�  �����g����������b�g��D���~��{ ����O�iD�! � !.3&.�(.&'� �%.b %�3.b ��. .&�{ !/3&/�(/&'� �%/b %�3/b ��/ .&�{ 2 ~"��l�!�~�&��� �,qb-!f���w�!�i��x!&���y�!�i��z!&���{�!�i��|!&���}�!�i��-�K,�/��� �-O��� �i,�K �L 3�,$���  ���@ ��MA      ���L �@  �N����"� L ������� ���'ݟ(Q������M�����S\W�f�3a�Zw U?���"� �� �� `    � � �� �               ���    ����M                        � �r ��K� �����pIfjqfr�bNSfYb�������1x�L�i�L sLb ���;yZE�L����&�"��;��E��/���b!���;��E��/���b��/�;��E�����,��s���� /�p�����p��ﲠ���p���y ��p��D� u (��|�/�>�����+�*� � 7*X�?�M��By�w6$5�*%�5*�s�/�9�&��*����Gt�"v�v�!uub!t⨤�u*)&5�*�4��w6w�'�w{���� 5"V�"��"�-#��3,�3��3��4��3�F4��D��D��D��DQ���r�Mb�����&��;�nq�r� x���1L����nM�j@      / �@ e�� ���"�1�q�Jr N�s��+�t�b �*C�$5�*C�%5�*C�&5�*B�+t��) *�C��"�uub��/���tub*B�+��&�*C�$*�C%�*C�&*�C$�*C�%*�C��ttb� ި*�Ct�� ި*�Ct�� ި*�B+�+��t6�&��&Bt�!��������*)B���$�+�?`��������g�)�v�vP.@@�v�Bv�u�tub *�C"�u�bvF�v/�tt!.u�/�u�*C�"u�u!.t�/�u�*B�v� ���+s��+�t�b�" �*C�&*�C&�5*�C$�*C�$5�*C�%*�C%�5*�B+�G���b'�  �*�Cs��+�'�&*�C$�*C�%*�B+�=��!�z�<"�i;)_� @� G����l�'�  �j*iB+�G'��&�� �*�B+�s�/+G��)&�  ��&�'�  ��'�j�/*B�+s�����&�'�)j��)؞'j��*�C��)�&5�*C�$5�*C�%5�*C�t"i *�B6�4���۲��/�����&����&��/�۲!����x������ �   ��T@� #��"�� B)�$��&��$�5*�C%�5*�C�����Gt�"v�v� uub!t⨠�u*)Ct�v?i���tub*C�>+��)�J ����Z&-���b[�h+�#��>$9þ��&���Jv&%5�*C��J �t&t!.[" *�B�� 8;�9;�*� �;D���� �:����z�'�+�����&�@���J �@� ���E.��J����Z-i�&�[&	&���"y	�z�[&�\&K[d\@N�J �P�[?�tt!.\�?���[v&\*9B��J�![���/�+���)�w��/+�+�����4���+��������+ �����i�KN�K��"�����+��d͊��� �� T�Wf��D��aI���J>61� �@  J�g0J��v6v)u�ju#I$��&���u�/�Ůtub*C�%*�Cw���/�w���/�t&"v�vu&w�"����v uub!t⨸�u*)C?���/���tub*B��t&�+��v&��uouvB#$���&Ϛ�nu�/�Ůtub*C�%*�C?��/��tub*B��t&�+��
Θ�� �M��8 ȿ�4@�02̢��Z�k��~�Z&�P�Y&T&0��R�b��{��H��+�H��+���+��(�����ǞZ�nPbYbT0i�^�R���'�H���v0i�>9,��+ž��"�Z&�ôv�bҚ"u�u!.t�/�u�*C�v$I��&Ӛ%5�*B��"�F�i�h�+Ii(g�**bf"&*e"B   ���w�aI�����f� L�H� �R$�5*�C&��"�u%i�u�*C�u� ��/���tub*C�u� uub���)$5�*C�&��"u�%��u*)Cu�������t&u*)Cv��tu� vtb!v���u*)B���/��&��*�/�/��&��&-3�0/�H<�e�J,֚+ �� �����K��� `!��k \� hH=�<��� � 
`�  ��xY��1x���w����V����&�@.HP��䑝��D.��+� � �uub7I��.��~�xy���M��;�d;ف�ޟn&En�D�wn&En�D
�E��D�Ev�D�Eu�D�Et�D�q�x���D�#x	���A��Mxȟ1I�����0�����&�����k !&�/����? ��� ���/@ -3�0���YrUfbe�/��Y�kH=�e�J,��30�/=�e�J,��+�x����?���

c(��w�/���kf�Z����	&	!.�l&�l�m�bZF����b��i]kb]k&]'	�J������"��*�3�̪�U�\�@�BA�C ��Z� P�����]]&]'	�J������ .M���L�X�b@�����nP2i.���&Qc&Qd&�& ���$���#��dO�x����d��Q�d�nZ!��cO�x����c��Y�UTbS�jR�J�c����������&!.�/�;��E�D		Ϛ1���/��&x�����}ܒ7;� x	�1��I��}i;��E��N&+ ����f�T�J� � ��F-�" �O�pJ�� �� ����+�r��j�~P2iQ^&.Q�_bf`afQc&Qd&�!����V��c���x�����c�jP�/���K(/��?�b�x�����迊;͝�;��;��x��1�Qc&_O�x����^�_�j�ϊ^�K�b�P�/���K(/��?�Y�UTbSRd���h�~�]&]�2���豲�����⮮c�����f�w� ����V��Qbd�b\�n ���K��$i�'�"[�[�"��nZJ\���![����(/a�O`xI�P���K�/�a��}����;͝�;���Ҡ��;՝�;��;������nZ�����;i�;��x�F����K�/�;����\n&En�D��Z�J�\?�nEn�D
�E[�K�K   h�`�} ���h�  �K��'�\L�d���x�����d�j�Z�J��?��x�����K�/������};���Ӡ��;��E��zK�/�;�E�KD	�
K(/��?�x��1��?�G����s̿d�G���6p�kLM�G�՚������ �:������l����כ@��� �   *��,�j��; �  �    �
G�� ��w������(/��&�Pn�.��b1��(�(O���� .���F.�� �       ���/��K�� �eeb!f樱�YU&�Z H
���&��&�Ƹ�ψ �$+�5ؘfe"����*Y.�f�e�/���Y�O�*���Yb!Y���Y!.�/��� ]:���]�,���1P�               �	�8 fe"���eD.�e&e!.fb!�e�/���fe"����e�e!.fYb!��(�Y�kfe"����e�e�e����f�eH.�f�e�/�e�Ee�e!.f�jY!.�/�f�eH.!��Y�k �� �����6G�� � �΀N�δ�a�t�b�t#)$��&��%�5*�B�������O�O@ �ƈ���� �R�f������P(/��O�ǮZ���B ������"H�������"ǀn�T&!.T�/�T�!����YD.�Tg&Y�'�F>�T��kr��3llsl!>m�{   �����"F���
.��&��+��!�������-���� ������ҁ���Ҁ� ����鸫 � }�	 EL�K���� �p@i ����F��6�O��n��b@H�J��b{(���z�&��"F����J|�J��/��|�f��&���F�� � �   L� (��J��&�	&	(?�t�t'�J��7��7��7��7��7������ ��B@���Ⓚ��(��������JX��    (���T���H��� ���c���|�E � �䀍�@����n��#��b�!.�h/�!���d�F)��J� ��:��G���4��c����I��� �
� �p����(���@/�F����&�Ū�Є�����������k����:��&,�p���p�Bo�L�"��"�����@���4F��!����y��
��@>��H��H  p�����ö����!��p����"��pI"���I�F&��j�/�'�"��Vwb��/���J J���Z�J��V� ��%����V� ����;�7I��D.�,  �   �IF6�� �I�K�I�Il������]%i ]��������J��d��*��h��������!�������SҶ;@ ����̠�Jrh�c��/�����/���9�&��%i "��W��29�&��%i "��Xx�����w7)M�J;��������K�/�����/�;��;فE�wD	�	�����/�;����Eh�D
���2�����2����;�D�;	D�;	��EV�D�EW�D������� ����� �M��1 �
�� N�K0�EX�D�͉�S�/�;����EU�D�ES�D#�͚���2���;���E�YD	(E	TD	-E	ZD		qr ��/�;� Mx�����A����?�x����W��(/���(����/(x��1��M���2���� � ���ϰ	DA�0��0,�� � @` �� 5N���@1�N�� 5�N ���F;���� �N��K+�J�J�-����J6�Z���JJ&J)��'��D�&�'��˚��J�nZ��J"JJb����rʁn'$��T�#$��Y�#��l�N&x����&�?i�JN�J����g�ZV J�
 ��V��d��B�+����b!�㚚&�	��R2C � ��A3�8N`!�R1�� �DM�P�ᦵ��� ��E�@� �݀��ރ��ۇ�K�݌�����ۑ�Kj�j�-�����9&���%��}S��'���߅tO�5A���	�P	�T �AN2�8D�R&C ���t�0R�MT R�	��	1�8VC`�@�u�HRM TR� H�Rq�HT ��  � A��� 1�D �� 1��D�   �ńs���T ćVC`�HN�QT�  ߁q XN 1�dă`�`@�� H �R�  XS� T� @��c] NT" ��=8 	� ` R�$= �S� `_ ��E@ҷA- ���T� � �N  ���  �ST�`R��DT�`R��D �� @� � 1� �MuC��	� @� 0��sLD= ��@ͷS�$�8 A� @ՅsCa QR�ՅsCa Q�1L	�� �S�$�8��C���N�Rנ3R@$�VqC`!����� A �`3�*�J ���b

�
k�,ْ},	� ������R��uw#&پ������&��!��"��          3>)�%P퀁� F����G�'�8"�b
�� F�������ho�����&� �F �������6��î�b��������� �����c  ��DO�#�8(�#S�`C��E`V��� �N$ �U`���� �� @�΃�CA��S�E.1  �B2���T� E�`P�P=h�@�