����  �?<> < |   '?
'>. "

	.       
 > *
0&0!*0"*
66'=8 61*62: .      &0(='; 
!%<>(+
;> +':'9='9=%'8'9=&'8'9=''8'9="('8':$?.!'7.!$?.!6%'5/%   ���(��bJJ�J�茀k  �   ��b���F.D����"� �    ��	6	 ?��������&�{  ����&��b

�
{��[�����[�� � �	� � �j��Wh�W͒k��� � m	����&��&� ���b����"��+ &!�����   �����"����pݧ�W> nb�@  [0�� 
 @ٔ�MA�� ���L�@    �ڶ����E!o�� 
 ? �� �� ��  �����|�� �    �                            ��_ ���"�*��������wŀs��r��s��O�2��"��" R�� �� �� � F39K3B=3'/3#3+33	3�ު����O�������������������>i ������������e�g�ee�ee������2�  ���㼱d��7��K    �������K �� �>�/�>��������������ݻ�� ��Z��4&4.��G�i�u�(��� ~� ���B�T�/E��e �T�6D�� e	g�en����������  ������(/�!���/����~��k�� (����b��{�����v�e�g��e��   A�2P N� 4n -�K ���e;SWn �� E�pJus �խHt�c�%\�� �AP�CrR� 0                  %��@�|��`�  ��	&31&��6�&;1�����y ��� � ��!.��/����'���&'&�&� ��K��M��<�2O�Ԩͩ�ԥ� ��'� ��<⨓��'<�K ��'='� ���� ��?���N͛ �?�/�K�aԛbK�aԛ堮��c��@��b���� /��@� �P? ?`��؇��ߩ�� ���&�&��( '!r�������'D&���� �!�歗c@������J!��!�筯"@◗K   ��? ����:�b��r�aya`�&�:��Ȩc����r��{ AB�C�D�ȋ ���4��c+(�@��

�
d��#0(���@/�&"d@���J�@x �=��!�z<�ice�Xb9�@� s	u��t��� ���$�d�� ���4��b��d������� �   ��✜d���� �Cd)Dd)� ��%��� �$(� ��%�$��� ���7}���� �	H?������ ����͋ 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� �� ��� ����� ���� ���� ���ۑ�K ��� ���� ��� ��� ��� ��� ��� ��� � �� �!�˽�K "�� %�ƴ� �&�� ������F�+0 ��cϛ@�
�

��# �c����@��&(@��� � �
��)��&�@���E��� 0on" y	{��v����'��S� �J�g� ��%�d���e�g՛e��01&�}�_����1�Jm���>�n� ��01&~���1�Jm���>�n�/��01&~��|_����|�Қ1�Jm���>�n�iʺ>nI{�/�1�n}��~���1��m���>nI/� �� ���J� ��w)  J
�
��(��
	�� n�0�1�byit}���~�_ߟ��}i��}�_��>�n�Ǣ�1�Jm��H^�lk�{���>�n�}��eg�e�La�`��a��;?f.2&.:&�m��ƫ� @�(���~3�iKM�2O�b��3�3Kia��π�:3&33B2�i�M��2���b3�Ka���cǛ����}�   �
邼����� (DLa�`��a���<v.3&?Ib2�b;�im���L�a`��a�����Ir2.b3?f�;&�m���� LYaN�`��a���?v<-b3Ib2?d�;&�m����La�N`��a��?���'?-B3Ib2�b;�im���B��݂�����6��I��h� �   ��)��9� ����������;!*bd(&!f?hg�	�� ��ѥ����La�`��a.�3?f�a�m����� ��2&��'�9&�;&�K�M��?�/b2���K��� �9O����2&�aY�L�aN�`��a��;?f-2&-:&?�Im�����La�N`��a�-3&??d�a�mѰ�'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[G�ʹ�����La�`ٜa��2-b3?f�a�m����� �&�'�=&�;&Ka��M�?�/b(��&r=Ki�M��?�b��2䒐���La�N`��a��2&?�b3?d�a�m��^j�i ������01&~��p �՚1�JmȚ�>�n�AҺP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6 4a���ίn���01&n�lp � ���n��no� ���n�#�bo� ��n�/�o�p� � �1��m��^�lk�>nIR�>�n����>nI�� ����������ݺ�݊��I�p���)�����Ŕ� ��/�� ����D����K      C �D ����R� � La�`ߜan�3�n4��ni1|481�J43D�m����/�P�� �� �� �� �� �� �� �� �� �� �� �  ��ڶ�ޱ���<������u��<�*>nI �C� ���w��r��r��r��{ ���"�n��"��b���# �@?�&2����+ �*�{��oyO;oRn� ^`��a�_]��b��L�a`��a�`�a���.r3?f��y�m����Lya`��a�`�a����r3?f��y?�Im���L�a`��a�`��a����r3?f��y?�Im���L�a`��a�`�a����r3?f��y?�Im���L�a`�Ca���'n1���3ai�3��_�����1�J�3��m��^�i��˸ 
ˣ 0M,ذ����[h<[, n	2n1����66c7Gb7761D����6��7�6��7��
33 0���44b�G���� J�"���� �J�"���� �{vJ�X��yI� �J�"���� �J�"���� �֚��{ܚ� � �u�t� e�g}�e� �� ���<��K�����d������v�}�s����geg�e�� �n�P���;&K��	H?��������'?�/�b�K�_����ޤ�����d��>nI �����'�a�_������J��&�J>�n� ����N�
.

���@����"!���`/�����)� �X              ��� �� �  0lc,�P��2�1L��0�?7���-��� �e�g)�e��}��2�i�(�(%})_���2�Jm���>�n� ���}��2&a_�8�����(�(ba�_8���2�Jm���>�n� ���}��2&c���1&�(�(c��_����1�J�2��m��ث >�n� պ �� �����������ߺ�TRN�!    ���N�R� �� �� c���}��2&���1�b��c��(_���1����2�Jm���>�n� ���}��2&a`�=��;-b3KiM��_����c�2�Jm���>�n� ���}��2&a`�8a���_�0��2��m��^�kj�>nI ��������7��                        88�pp����#l���� c��eg��e�eg�e���eg�#e�e�gi�eY���eg�^e�e�g7�eY����e�g �e�eg�ie�Y��}_����e�g^�e�eg�7e�Y��Ūeg� e�������})_���}�_��ٚeg�^e���}_�����eg� e�e�gE�eY��}�_����eg�^e���b���� ��� eg�Re�Y_������eg� e������ee�g�e�L���������'�������!.�`/��N�!.3�jYW��X��U��J���z�?����??d���e��;Ki�M��{��v�JVi��z���d)�d)e��X��ȣ� ��/�K�aޛbK�aޛ    TT Q��PYÐ������ � ��  ,- /�w�|(_v*�w(��*�X�*ubtb"c!*⨡�"�J�/vs��"�rq)w|�p(�"(?o$��n�n�&!'&!,2���w�Po�m���hÂl}@���lt�$$bp ��X.��/!�x!����"k0�!'$�J'j;P"F�i�h�+Ii(g�**bf"&*e"!*bd(&!�;�ӛ�����T��؈	�CD��@�������%!.cq9|&R!q�|o[  �%�&-bp(�b)�w$����b�I�H��AG�q? ��lI��4���G΃��R0 N %�G΃��TT "��" ���b�I�(H��	 � 5NT"	���N�B@��"mI��4(��GL #� 5�)E �"mI��4(��GR0D�#��"�S	�EE) ��b�I�(H��b�D(�8R0	���N�B@��bmI��4(��bmD�ԃT�	���N�B@��	��R�H�RDmR���@��@O %�T�	C��4�DI�3S� s\���R�R�N�@p ��R�R�N�@0���K�D	�3 0���K�D	�3  �N%�	EI�3S� P >�R C�DN %�T��A�T@΃�S���@RS �S� Q5S� 	S�8E �ES� 	S�8E �ER�C��`� 	��4�DI�3@N���Ca QN%�PE �SՅ-ORQ��5` N���N N�TP U��0� A�Q`RQ�4N %�T � RC �TNB U� @����DN"%S� �T�0"��CS���D�0O�#�TBȠN(�U�$5�`%6 ��RB 4N %ER��T �C`�T ��4N	%�8�$�RS� Q� 0 � �N`!NB�T΃�S���SBRS �R C�CA(S-O��E��IA�3L	�R1��SO�#�T �1hI �	�� 	Q � �PA��G S��C��U �#�N�@�O�5N�P��R1P�R D0N�P��R1P�R �1�I� 1�8�1@�S��C��U �#�	� 0P����� D �� �����;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    ��}�tq�on�m{�| ���������������g�ݛ�ܖ��y��{~ِܠ/����&��I������   � >��y����� ����� �	������� ��A���D@��
	�gh� f �Š/�Ť��7��7� �����/�������)��)��Y����b��i��F��6J� �!�⨾���2Ⱥ���2�����0��{��)���� � �� �D= ��@ͷS�$�8 A� @ՅsCa QR�ՅsCa Q�1L	�� �S�$�8���HP���	� 
� ��R�� ђ���y���Ҵ` � F����&�� ��)�.�暎J� �   ������ ����)��J��   �|�A�|����Ũ�� ��� �� ��/�� �������'��; �� ��� ����b��y�N�¼�F�K��O�F=3$3 91��	���� Agh�f���� ���� O �	��I�����b� �   ��b����&,!��"�ʟ�-� ���ڲ�ދ �   �l�Ao��n��&� �����?����Q��Y���)�\���)�_���)�b���)��� ����ȟ�����y��C0 ��LD!  ��N C�� �Q�> ���������J��I&׽*h>F3�>d�M�����R��� ���� �� �����;��A����b��c(����?�����J��?��������K��C�����'��"��c��k    �
�}�tq�on�m{�| ����ʪ�ժ� ���y�������g�����y��{���������d���� � � ������� >�{��X�g��M�ӻ@� ���KL� J