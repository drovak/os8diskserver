����  � 0000  . A( <A-0
0728 8 8  -=��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                     _ U��MA�� ���L �         � ��@  �   l ��? �?p ��8 ?�7   �/ ��  � �� �� �� �� �� �� ˨ ө  �������      9"��� 6���      � "]Z#֩A�?���s�
���  � �Y?����?���R��`  ���

c��b

�
�菐(� � � (���@/������ ����*� /������&!̥���"�
�?�������  � �6� ���
�)0�c(��'0�c ��J.��
���&��H�'�.����&��H�'X�&��K      0�� u (��|u |)�ظ� �� �(?�r�� ,
���,f�m��� ���"b!⨘��*��(�2&/&"��(?�&�!�ʠ������- b'" �&��-�-�E� .(Ҁ� �--b��� .&(Ҁ� &F'*G'�- ��I�F$rGr� ��I�F'"G'�- ��JI���F*rGr� ��I�R �         �,�!.��!.(/���#"Vk��-"-b ����"Vk&-Vk $b	KbD�%K&K	'�J� ��-⍀ޱ����ڒ�ډ�� ˀ�O�m N��ډ��P � �]$b"b	bcM	cLMb!L����J섯#���! O�j]�J�#�(���]� ^��Q����؇��� �Zn\!l�"�����,�j�)� ]�]�J��� HK`��\.Z,  �T-�-."TO�12"TN�56"Sc�0X0�`00Ƞ0L0 �� �T-�MN"TO�QR"TM�UV"TL�YZ"Sc�0X0��00� 00� 00 ��S�cN��	��� � ��l�Ub!�l!t=��!�z�<"�i;)�f��H/ T	-��T)]��S)c�`00 �R���D�0�0 ��²v���q��}�� �':"ȇ�q�9�/���{z$�8��)�7��6)q��5&����9�/�8�I�� & 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� 71�