���� � ��'=%(7-	  8!1<;>(*+'2	'8 (2(<*+
1>(*#	!*.  <;>(*<	!*7.1  $> +8%>(/%
%  /u;6?93&v �B ���������                                                                                                                                                                                                      �'�B��t��s�������e�
�����&��� 0�D��L�LI� �I �kp���F�D.�&��(���c����(�/�S�
U)q	w�7�(S
�U�qb��q���{�rw�l)��AIkl	�Z��[��!�� �����x�?������e� �x���>�� �x��F������ ��� @Ok��(6�(B(("&&Tb��_9]��Zym �I�0/f����0�/�h����/�0����0��/����֮�Ɗ@Ik D��&Tb��_9]T� ��_I]���N� �A� ׉� P�O� �O P�ք��8�����ELc� I`��@.w�/�I�KM�Qe�I��m���q�n����vrg�ǁ0�/����0��/��������{��ĸF ����8�Qa�I �A�/�A�S\�]��K@��L� �IL�S �I��BIk $^���_I^�� _�]���p���Y��P�&F.D.�"׉l��6Q �B�/I�l��A�Sw�U�!.$b!%��L@�w�/�<��IW�Ќ1@ �|�!����A��b�&�B�.XiT��)�&)�Bh]�)z)qq�v"�c�+r)TL�))$h]�q��OQ9q�
�'Tw�)h)]q�w�qw��scdl)�Q�#��Aqiw��Sw�U�(OIQ���Q �� �B�/�B�qL��)�)zIqq����z]��A&.Xi&� � T	�s_���� `������   �``�8�n&A.bw�/���Zၨϳ8�i)�a09c(���lT��fr)N)+r)�r)]9����)h)�+rr0�������w2Y�H���Q�#8��I�T��))$z��r,�r]�I�H���Q� ��
�(��!. /�������٫�ۚ�W�T])ZM��\�+r)X$�IR���A@�(D�����ܱ�d�c!(�D�B��l6�S� U	(�S�z]9QF�QI�T
��r�c�]T�d"_��D�<N]�Tw��_)]Q�#�� �ødH.�g�g"&S �8�/�9����^��c��r)!.os�+r)�r)]��U����r^��_)]���S�k�� �L{� �L�� ����؀� ��� �.��}�
B�Q�I�`��f����Q��Q�7I� !��b�bc���&'6�'� (�(����2����a&�J� ��b�bc���'a"d��� ���d�$2����.c%�/�S�
U) �M��`6	I3 �UL`!��CN�!�          S	PRQ�	A� 0C���^�sf3                                                                                                                                                                                                