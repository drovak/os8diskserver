����  @   	   ! 	 '  	   	    	    	  !  	?   	 	    	 3  ���������                                                                                                                                                                                                             D R�v&xş��C ���G � �      ���  ���$�U` P    �            ���8 �t�C ���0���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s�
��� �v���؇?����� �����&�R�������k ��'� ��̕�6��C

�
�萦8��I��� � (���H/��"��� ���ú�d�/�� 	� �����}�����'����2���� 	������ڽ������!��� 
.

������ z (��~z ~)���R?�N�@�?X��U ���ė��y��������z�& �&��&��     ���#�b��&��Á����?����z���
�l�
'�
'�
�  � ������� ��/�����̚��K�k ���/�!��� ���/���ش� ��Xp@��u@ee�q�}��	ȰD�D�!�����?��� #	 4�
����@�␠���rc����"�j����/��	��l��[�������� �	����k ���4(���i 	��5��K����iT�� �'%f(?�&�&�"@����'�/����{%D.%%bDD�%%&&� %'$�%���K� /��@� ��P���9  qJ@  �	�����m��������a����������!�����ǁ�#�=�J�]���à����'��������������s���Ƞ�� �������	�!�̘��ډ�������ǁ��4�������y<������ʉ���yN����փ�����1	ɑϽ@� 6���������;�����������)�������è���& �����?������?��"�i�������è���<�%&%�6c� ��������2� ��ț�) &�)�����4(���/�פ�ף  ku�D� ��G	F��E �?��*�� ���I@AD9�@I������������!>�����Ú�����I�� ���n��f��&¨&��@���/�O���ʨ/�Ȣ��b�@/��ʨd˧J��/�Ȳ����/������      �h�u���b�#i� 
(���J����J ����y� �((b

�
�()���S���H�O	�d )��@1 ���ǁ���ş��X���������|c��i�q�v�{���������������!����|����������|ę��������w�|� ���!��&��?�ܿ?�>?۾?�=?ڽ?� 0��º��D�� ��J��%%c� �H�K�����K  ����IH�GF�EɑϽ@  dD� 
��6��L
�t���� � �	��(�����0�ۙ���%�b&c(���%ǁ%�&�J�&�� �/�"� "D"�P�����<��B�\�;�������ǁ���/��������i�������������������&9� �
(�?0��M`3���5Dɑ ?Y���@ϔ> � �	��)��y�������p���b�j��(��(��(����� �s��¨��D������ǁ�� ����)�����7�������3�|#�� @�� #	� ��� ����&� ��%��'6ՉL%�< �%'D�ի~,�(/��kr����$t	���ID��f����	� � � !"�b

c ��"�/��	I
��"&"D."�"�i�iC����� �����  "f�*&�+�)c�(/����((b�(/���@�����("P����)�"���)H.*%&(� ���%�%)t�+��*��*)�/��K �
!��&����&�����J���� �? ���?���R��`��@�� �$��&���,l�k��s_�_�_�_�e_�v_�_�q_�}_� ��r��/���"���w� �$�J�)$b���)�"���C�������h����/���$I�$�%&%9��$����� ���4(���/�ݤ�ݣ%%k��&(?���ؾ�� @� �A����� �����s��|����������� ����^�&�&7�"Ț��#� 4�
����@������rc����"�j����/��	��l���&�&7�"�������k2�J&b�bbb�j!.�/�a�d����w����w��r  qJ@ ���D���J	�K���    \ P�@�����  P             P 0         n �P 0                              �ӛT���D�م���������������������������;�<=�>�	H�IцE�C�DÐ�Ż �� @� @ ` 5   @�D � � @p q  r s  t u  v w  p0 q  r0 s  t0 u  v0 w  �p@ �q  �r@ �s  ��@ ��  ��@ ��  �p@ �q  ��@ ��    �    P � 0�p  � q  �   Tp  Tq0 � ��L � ��AL �B ��CL �	������{v�qi�� 5�E3��@N$ TA���ŠTE�d�8�1ՃN� R�?E�d� 0SR���MԄB	�SA�RM TR��  �8C��MAx�L`!ԕD�RDVCS N$ SRA��G�LRP΃T�#N�`�N��A��PM�@�D	�T5 ��PԃL�`���@RDQ 	��@�`6��0	SAR�MTR�0 ��PS�R�MTR�0 ՃS� %M� TB��3�RA��D�D@N�!���1(v(��D�_ �L `� �N2E�_	���`�e8`��DA �N�HVC`�5�O��HVCSV``�N�HN� N �RAS���`Q�6E��OB�N5�4ՃV�``��3�N@�V�Cn! �N�HVCS��N �N�S���,��,��5 ���N� *CML@
�L@ `2S`Q�N@�U�S N ��dR�MTR� ���HUS@"(�"8��d��`��3N�!R`�	5��4  �"8��d�L��5  �3"фA�T��S�L� ��"фA�T����C �N�	H��C8L��AE� K�8R��R��8�3D��U�S"��`�3�$���3D��U�S"��Y�4�?S(S�`SSAN? ��MA	:�  �=N�S��D  �}�� � ����;  �����  =��SmS/��  �}��� �  �T���;  ��U�o2  � =�U3��; ���OB��3BR1(S���@TDT� �$�MA��{	n123��� ���TO�#�CS`�(E��}�l����T�`
 SR�GB� 1��Mz  �`QSRQӄG�# �E	8�`@�1� �E3ń �T���4 T�	����@MN1 TP	���CE 0�υ���@RM`�R@	�ST� N �  	X�R5`NQE%��4� ��SE	8  `Q�SE	8 S��X`� ��DN!	�Q�	� 0�D�S1��nhC�ML M��� 0�v ���DV`!�0 5`ÉDVB`� A`6��8NR�� P��r���R C�H�U3P28NS! TS� �PR�I�3 Q�U��j��;@���3D```��A�!T�R�S O�H�#r ��R �NB E`��NBTO��1�DA L  �1��D�"8�AEȠHL� QR���C� �S`Q�N@���H��8�T������A���DT�0(��A) 8�8Se`4SN U`�hRM TR	��SDQ҃"����HXTRI�3 �R`����AG�N�$�N@�	����Ѡ�C��4�MAV�CS! v�҃S�`S���MM3a� %�L��@RQ@Ä�E ` 	58�5`��� �MM3Ma3@���N �	�$� �AA�H��5�l@ ��8 �ՃS� %  z�C@@ ���0VL!`a�  �N %T�/�UDN	L�M5S(`�c� ON U��5�SE ;NQP�`` A���X��0``��P ��a O`�Q��C̓T	��;NP�@(�E�O�`�SD�4S�`�T�  O`QMa6	�N�	��VRT	b� 0`Q��E����E���D �hM`!� #@�`G`I� Ό1C%T�   D RR��38  � �� `� TR��� Z�	^���� ^�� �  	� ������£�                                                                                                                                                                                                