����  � @�                                       $*  *$                                                                                 ? ? ? ? ? ? ? ? = >>; 8 >>= A18! = ?8?                                                                                                                                                                                                    3�    M �      ' �         � �� �� � �
               �4 �                      � Mc       X  U            �                                      �s�
��� �!@���? d����:���&}�j�?�ieffy|�i�I?�/�}��e ��}n��*�wF�giwgg�b

d
(?�g����
6e��f�����������������}��f¨�����ORf�&�����S(/��TnSMiTS&M���cI�cH�c0�c1;i���?�)��|� KV�����z�ǿ ��JЫę� �[\fJKf�7b�i@�&Fhb���{{�74&4v $4b
�v#�˒H���h����.&��(��4n_4bv$4
.v�#4c�u�(���(/���(���(/���(���(/��   �H.�H.![�F[&hFb����(/KJF�y�|���J � H�
�
������ � K�����������/�3��$��2c3#b%$b&%b2x)�%�3&"���4�9��/�'RE��G�?X(�G���������   F�Nh�/�'�{(�{�� x	�&��G�����и��K�t��b�j����b�j����b�j �Gw '4bwF�''&� �bbt�ݛ �b@/b�b�; a a�a�i� �a�Oa���Y�/Q #&J�� t�&(#bx9�%�$#���4�9��/�'��G�n���@�/�\��'�E��G�?�(�(�i�䄀� �($b&#b���#)"����(�%�) ��#"%n$&&&t ������$H/�&����� �����   �  � ��  �����������=��!�z&���1@�T6 ^�1 �(b��c������-v0�-'��t->Ƚ��9��/���--7������C���C����@����C����@����� �'&�->���t v&�9��/�ڮ--7�������"�h�H� �'&(�I������ ����@����‾��)�&�aQ"��8��K ` � �D8� %F�&s"G�k � ��_�9� (��J�s4&4�&�4rJ�vF�(4b�(G�b(4d4v ���4�8u�/���'D)���4��4&�v ���4�8u�/���'D)��u�(̋{   �s�ib���i�b�b�bc ���Jw�H�������5&'������6&'�� ����������� �(.���%"x���(�r(&�(��(��(����J(�'w F�((&� ��G��������(�'E)���� �%&�G�����'�E��������!.!@/!�(�����۴ !."@/!�(�����۴����K� � ��b&� ����a�k a!b����&}��`�$��A �
� �߶D� �1��!!�@!� ���� !."@/! ������ �!.!D.���!�"b! �D���!��cb&!.�/�������K �!.!@/!� !."H/!⠸����� ���!!��� !."�/˔���K��������������������� ���&�yÉ
Θ���}�   �
邼}I��@߶D ����@AfBbv"J.v�!b!x)���"�x��J�.s�c������@CAbB�b�����J���    �/0&00C(����b!⨶���9��/���v �
.v��c���(���(/���(���(/�������@���/���@�/�!A�������A�bB�j!�;Z@O |A��?`�Od�@  ���?�_�H�����_7b4b�rJ�v!v "4bJ�v4v  �i������_�ɶ(7&���@�(�������?[�K ��C)�67�{ ��C)7�'� �   �)�=���~5b7�b.�b/�b-:i� ���=q��6r7�b)�b.�b/�b-:i�� \��l,�+�	� ��K8D�KA q�'���/&��� ��'���/&��� �i�I0)0C)1�/���!>�>cw+),)9)19&1v (����&������"��"c!>�>c��/!�>2>�jt b�&7sH,��+������*t bvc!>�>g�?� ?��� ������no ���	� �i�H91&~9�~,�~+�1�/~�~0�0C)(?�'>">1bv(����o���ƪ����!>>>&�?�u"s>>&����"cw�����*v btc!�>2>�h? .?�k J.

�wsbws�k �Rt"@��v�+ �>&�!��/���W���f��@�
 !��bL�/�����L@/���ȗ��L�H����/��D���   ����bc�J>>b� � �	�0`�i���>`"�`��`�``b�L�N�)�Ċ�Ī���`�+�)`�+ �]�/�h�F)[)�[��hd��![���~[�~F���+[(/]!.^!.�ț �B6� � �gK]U߀	36��Έ��?�� ��)R�NR�/�?����q�'[]f^cfN)ON&�9F)`)F]b^�][b^[fb)a)R.���q�'R!.S�/����O��J����K�/���z1�z(��0�0I&1H&���;M�<�� ��z�z���ϫ �?�/�?������mF��B@���Pn�����彀]EK�W݀� S�)�3�94�7ߏ���P�)O�)P�)LOb������PO&�)�0�
1r
�~O�)LNb�������R�����������d j �jd�                                                  �RD.�
&ҷ�������������`����� ��`��	��J�g�v���V��>W ��O�p�3h�⪀O�P�j���P����RR&NO&~!�a /~�!b� �^[&]^&~]�~`�~F�~��~N�~����)R�"�P�zz�� �!��  ���=?����6�)�5��@�����)ccB!d� �c�)�P�� ����� ?�����&e�gg�gg�gg�g�������
�y�¹Ҁy�݋fKa��fͣ�3�u� X��  �	
!>Fb!��(��bDb�c(��/��D���b�"cr!�D
67
'� ������h!`�`qb��b�`�`�k �ft&?�(/�B���JD.D�� ��&��&(������"``&�D���[�\c�d ��+����`"`,b��t`"`�k  ��?���?8� ���g �=ɓ(�������)A�&@(/�̶B�&��)�ɢ�A�!��B�&@(/�̶��)A!.A�b!@����@H.��������9A�"���A�"��A�"�ɓ!�����ʒ@��!�� �    �	=s���b��b�(����������D��� � ^���P 0�^F�P�C  �^F����  �^F���ݺ����Ê�U �?�/�q"��f�=i��(��&����(O�����8��/����(������B!���������cwF���cw�j���H��F�!�迀+ � �       ��&�&�&7�J�&�&t�9�+,f>�k�S�����'��J������ ��.��qߧ�� O���?�I�K � 
�����n�l�(����b���)�"���O���(/���(����/���rH���  � �&i���� �	$����ˀ��!⨱��)���j�}���鱰����|���{�����5�s���ܩ���   �C�T @�LMT@OReփ �S�$�'j�s`��   ����F
>

����� �w(�u�H���)� �&!̛"���� ��)����� ��b�bl� ���b�(/�������+ ������)H/!��� ���&.�v �)�J� ����ݛ �R(/!��}i ���� U3�.������S��'��� �@  �IHf�����F�������J.
�������(����F.����/� ���(���(/���(���(/������H�j��/����/����Ii� /��II&�z�1zi(��!I���I0&H�/�1�v!H�/�;�|𙀀K IIi��� ���3�KOI;@&+OVw��81���/C�O��?�� ���&��&Hv ��&����������"��&��&�I�

�
��H�/��"I�������� ��v �)�
.v��)���})� �    �H��t�/��N�+ �H��t�/ƀN�+ �	�F����J�/��"}���� >��{? .?9f������d�OVw?O�g���� � � �����  �  � �   (����b����������ߒ�������� �   ��ZtbVZb
tbW�j�)Y
c(��HY�H!�u(/���(���(/���(���(/��������"��"��"�X&Y�/��"X��

.v�
.����X&X)X)W�JZ�tZ&V�J���@1ê�� ���� �@��������w 	�Z&tV&Z
&�)�W&�*�(������!.Y�h
Yt����(/�������Y����(/���(���(/���(���(/��(���/�ժ��"��"��"Y!N
�zW�JZt"ZVd�,�+9f��뀛������ �W�K׮� � A��8N� 1��a@��ʼ����� 0��>P�����w                                                                                                �d j �jd�                                                             ������������`����� ��`�                                                                                                                                                                                                