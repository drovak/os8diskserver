����    @C0 ?<h   0	0=
; 
 ?>(**>> *%%4%1(4%1(<%3%1(?	%3%1)
%3%1)%3%4%.?*1%8*1%.?. ='</'<0. 
- 	    :   :   :   : ????????  %4%1)%4%2; /	 �� �������������������������K ����� .��d��J��d� �    	B1 �� H �� ��/�� �������'��; ���6��C�(�@��

�
����0(���@/��"�۔� �   ����� ���&��'����@R��R C��@�?����� /�! �w����          �          <� � BlU�� � y�w|�     ? @�  I� 4UjU� h$������������b�                      L VNP   ��"�#�<^Q_ r`;r => ?T>/=,�l�a�<?+@ 3<��E�.������ ���bL��D��{(�w� �(w� �w@�wH�w�w��(�w�  � w�Hw�@�w@� � w�w��w@��w�w�w� �w����w �w� ��w� w� �w �w � �w�(w� ��(�w�(�w�(�w�
(�w�(�w� :�(w�w�! /w�w!�:(/w� (/w�::"w� � w�..". . w�w�44"4.  �w�w �:(w�:  (�w:�: (�w.�4 w �!(/w��"(/w��#(/w��$(/w��%(/w��&(/w��((/w ��)�(w��*�(w��Y�(w��-�(w��1�(w� ��.@.�w� 4� w�...(w�4.w� .� w�4.4 w@�2
.w� +� w� 2�
6� w�+.w� 2� w�+.0 w@�'.w�( /w7��w �( /w �:/ w�Q � w� Q� w�./Q �. w �./Q4� w�@ �A�w�  �wQ�(w�Q ��� w�w�Q �w �� �w�w �Q �w�:J& w�w�J . w� J�J /wJ� w�w�J:" w�:J&JwIw�J /w��V�4 /w:��o �  �w�� :�o �w��w�4� U� w�K42 w�:M'N . w�MwY.N& :�M5 w��?L4 w�:�'N�N . w��wYN�.N&:�!N�5 /w �.&5" w�N.bOMbc5 /w ��J&��!J� w�c�� w�J& �J /w �@�@�w�Hw����
�F� 1�F,��w���� w�w� ��(�w �w� � w� �w� � �w�)�(w���F���w� w����w ��]� �jwɘw �� .P� w��w���)w֒ � �Q /w �No�N� �N7"@T��N���&9&� �DEfI.�H�QG� DA n��CQoB nJ n n nO n n nRc�� �� �� �O� �� �� ��J N�I���HQ/G$����@O� �J�!$D�SJ�����@�EOD �ED�EFE(/D�N$�S�@O��O O��O�תDD����S��JAS�Aob�SJ��C"Jb �A /Qob �B /Db����Rw9�H�QI���Gw)R�(���R�w��./Jw)�C���B/Aw)���G� H�IRc��R�)(䀾R80R�{ ���./�G�
.�R���Hb
���I�k��"� .*  ��m���
� ��w)  J
�
��(��H����%��d��������d�j�|�J��P��y���C������?���1n���?�1�v��9C����1x�<C��0�!C�(����ȟ,��<(I����D�Q�/��"�Qf��)����1���,񙼀�VyF;y���k\{B�����'��6��K{�/���{f��nGf BR ��<@�@�� ��3�� ���&��"�r&��'�@�.����&�&�&P� w� e��b�w�a � w� e�f� w�a � w� e�-g,.f,4b,  �w �e.�f��g4�b5�(��ww� e��&�,)bf`�w�Y��w� e���)bf`�Kw9�&<4" w��� �c��/��K���t �Tɴ��)�V ���b)bf`��w� e���)bf`�Aw	�&��  /w �e(�f`̂ �e(�f�` � a�w� ��JelJwIdw�w� ��f,`���ߨw� ���b�b)bf`�w�  /w��f)�f`�Owڒl e�./�g,`5�a.� w� e�./�g,4`,a5� w��$�&� N����J9b neP��g,`J�a7�� /w �JD� ��g,./�`�a �w �ze��&�&Yg,)f,`b�w<� w��& ,� /w �e���bg��)bf`�bw�"  �< /wȒ b�� w� |�e���bg��)bf`�bw� <b w��& ,� /w �e��bg��)bf`�bwɀ*�8 V߿Y��Y��< /w�� b�� w� e��&�&�f,`���w�w���& ,� /w �e���b�b��bf`� ��ww��& ,� /w �e(�g�΁,�c`� a�  �w,�gc�` �, > w�)g,4,'c`� ,�� /w �e.���~f(�gc�` �a5� w�g��c`̠ � w����WP��<|���i.�ik�e�52 w� e�*f,�,�c`��J�J�J, ?w �e(�g.�,c|` �#f,!g,�J&�&Jt�c�` ι&�J&52 w�J�J e�J�J
@dw�d�w� e�.�,(rg�fc�` �,a|5 /w)�f�g���bcl` �,w9<(/w5� w��& ���e��,�r�b�bg)�fc�`,�w���  w޶< /w��Fb�� �*� /w �e-�f`��� w� e�f�`� �1a@w��w@�w�w�Hw��wH�w�w�Hw��wH�w��w� e�`�a�Hw��w�@�w�w��w���U���4��b��n\����9ib�{d�~��"F���
.��&��+��!�<�9y������@������ �@w���w �e��f�`
�F .��a)��w� e�f�`�)�a$��w�a(� w� e�).f��n`�� ��laY��w� e��&�f,�&` �� �w b�� w�@mi���? ���s��e�/� H �Q��?��"[�"��e�/� H d�/�ôß�.M�^@��; !�@N Â��O�x �����n����������tIq,��s)tn���x��� ���/��� �檨D�����K    � 
��` �D  ��y� �Ȍ��+ ������s� ������d��0(��@�
�

�v���(���@���v)��J    �� ��� ����b��{kp&����� ���@�?����  �� �����;��A����b��c(����?�����J��?���v��vt���K��C�����'��"��c��k    ��}�tq�on�m{�| ����Ɉ�Ԉ� ���y������y�����gt�Ӏ��/����&�oI�p����   � >��y��� ������ �ag���ә@� ���JK� I��������6�rI��h� �   �v)�v9� ����������; �� ���q)�o��p�����TN"�  �� ����/��qi�s)�v)�uY����b�ui��F��6��J� �!������2�����2�����0��{�v)t��t疮 � �` �𱛚�U� HP���� �� �IK�J��ހ F����&�� �v)�.�撆J� �   ���v�� ���v)��J��   �|�A�|�����o��p� ����� o	�pI�v���b� �   ��b����&,!��"��Ҷ-Ա�̲����    y	 ��D�b���1 �Ei���6������� ��{��]�\Y� y@� �JK�I���� � �l�Ao��n��&� �����?�t�q4�q<��s)q?��s)qB��s)qE��s)tn�ȱ�x��nȟ�����y�����
��` �LD  �� �C� Q�� 茀������ t	qT�tr����AN2�p-�
��@ 1�o�/�;�mn 1��l":1���k:)����<�=<ݺ�J?� �a �   D�� p��t� ����Dh�����K   ��b
�I��I��   ���A�� ��A)��J����  ��b�!D�⭭4� �D'��2� p��t��K ^A^�A  ��� 9�@����&��"(����/�M����Aɓ�(O�@���������cɭbɀ���J����@/�ȢH��� �� v��.�xB�