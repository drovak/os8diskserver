����    �    }=B ;/��������������������������������������������������������������������������������                                                                                          ��נ�����ō����É����Ġ�����Π����Ҡ��Š����Ԡ�����ˠ�Ӡ����č����Ӡ������ˍ����Ӡ�����Š�������Š��Š���ō����Ġ����ԉ���נ����٠����Ԡ����̠�Ҡ������̍��������������Ӡ��Š���Ǡ�Π����˿������8�   �����mE���  0֭A   � �� � î "3?"��!!� �D�T  ֔A��8 0֔A���F ֔A��PP֔A�����֔A���� 0֔A�	�1 L֔A��σD֔A��T֔A�C�	 D֔A���P 0֔A���֔A�B��A�|A��T�DK���M T��E����� �	�������������Iҳ���É�Ɂ�É��Ҡ������������ ����� .��d��J��d�U�   < � 	��@�� H �� ���É�ό��ȁ���<� �������'��; ���6��C�(�@��

�
����0(���@/��"��� � � @�?����  ��! �2 H ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}on�m{�|q� @DLZ�]��g�ٛ�ؖ��y�|ˀ�ؠ/����&��I������   ��������� ���������y�����y������������@�����"AB3H@3��������6��H��h� �   ��)��9��� ��?�>��� �������C���������� �	���/������,�<�����Ҙ��<�|��&�Ҙ��ÉF����ǉ���� !�/�����/�����/���������k   `�H �P�����  � H��H@B3A�2��"� ��)����@O��y�����撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�f���� � 5R��C�;�~� �	�� ����/������  F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��Ӷ-� ���ڲ�޿ � LD  �� �C� Q�� 茀����������   �� �    ��HAB3@�0�� � ���)��)��)��)� ���b��b��b� ���'��B���������&���� �!�澣c@������J!��!���"@�⣣K          �������TN"�  ���㉨���K �	 ��� ����� ����� ��� �֔A���֔A�B��A�|A��T���  �
�8�2 �	����������� R֔A���� 4֔A����@F������@�EE�����@�������@�mE���  ֔A��� 1�mE��� P�EE����@F�Q����@D������ 0�  ���C�3�%���C�3��F���vr� P���wr� P� ���@� @� ��Y�B? < Z~�O��Z�� ��� p   ��1:" � ���/�  ��YPU3L  ��1�QTX]b����M��T� � U�w� C�\$�<� �vV�F�8gU�r      ���� ��������
�< �   �� �            ���    ����M���� �� �             �           ���{�i,����'�ov{AfvKbFUf[�nE�n]D��$��#�����?�@�G�i,��(��'�Av���KF&+S�dMb�����dO�����d�0!�X� �'�(��2�������2���!.��?���1ݛ��gh&Ii&Lk&Ll&mnf�&r�/����/���;R� [����D� L�� ��I��Z/>�H1	���,�\i�����b������"����/���b!�����/���b��/�������!.�/����\ J
�
����n\H|�c��k���������Q���T����X���b�]���&��*b���m��KF&�u��F�⠾��+����u�I��H�L���>M�/��&��*�/�/��&��&.+�*��?3�e�J7���.�+���[rW�k�?�4e��(��.�+*��4�e�J7�����\� (����/�վ[|��KF&����&�?u�JF�J����j�\X B  1�e1)�Y�� �1ś��L� �������������4 ��@�8�Q? �43� �#��c��k��!�"\F���b�xf�|����	&	
&��'��'��
!.	 /�[��H����V�*	. ��xe.~�j��x�~�j�~�x~"x	d �������"��"΀.3�<�U�N�)�9�\\���|���&1]�� �@_���2�����I�Cp-	ᘭ@�
�i1 jba0��U[[d�� .qpw��.R-i)���&Sc&Sd&������"��~�!��dO�����d�0!�Sd&�|����cO�����c��[�WVbU�cD���0���T�J�c����������i�����1 �ȟ,�0�Sc&�D>��)_O�����^�_�k��^�J����'�� �4Q3C�� �+m��9?�Ԁ�* �>R-iS^&)S�_bf`afSc&Sd&����X��c��������c0i��R�/���C(/��?�b���������1?��1�C1�c��,��b�R�/���C(/��?�[�WVbU�cD���0����S�!_�(��S�/�0���R�/�a����_a&0��b����_b&0��0�T􄀫8�iC��� A��#��0����X��Sbd�i�����C�f�"��%� ��"��n|J~/P!�/��(a��`���R�/�C����a�/����1�?��1C��/�1�G��1M�1Q���&�|�����&1X�1^�������C����1�
!.	:)8��|�J~�P�y9iy8	
9	C� � 1	U�K�w)K B[X��H  $B�%��d��������d�j�|�J��P��y���C������?���1n���?�1�v��9C����1x�<C��0�!C�(����ȟ,��<(I����D�Q�/��"�Qf��)����1���,񙼀�VyF;y���k\{B�����'��6��K{�/���{f��nGf BR ��<@�@�� ��3����B}�f�(/��&�Pn�.��b���(�(O���� .���F.�怽���"������1��1e���@�/�1��,�1��@&I� �  �    �� .����"���1��<��1����/���2��T�ne�b����ٴ1����/�1�o�+1��+<��(I�٫��N�6�2������ӻ����;�K�F �0�<� �S�F��6����QB �eeb!f��[W&�\ H
���&��&�*�*8UA�U؀U�Q��'��'���[�c��c��j��!fe"����*[.�f�e�/���[�H[&!.[�/�[�!����8�;	<=�o�/�8�;	rs 1�Oq":1�O�p:)�շ�6C �1	ȑ @��dqwp�r8�fe"����e�e�eਡ��f�eH.�f�e�/�e�Ee�e!.f�j[!.�/�f�eH.!��[�k�o�^h��g�hid�I�ivb���wO�k��L�kld�L�l�b���fe"���eD.�e&e!.fb!�e�/���fe"����e�e!.f[b!��(�[�k�Mq�`1	G��4C(S�"@Q8AU�	m �Ju b �T�f���]�R(/]�O]�N|��]�]�B ]����"H�������"��n�V&!.V�/�V�!����[D.�Vj&� �`�/�_�`0i��N�Tυ��@` H1i�9�\��/����/ݠ��/����/�1�->�1	1>�1	5>�1	:>�� ������<^_f;p"���i�����5i��c��F��6��/�H��n��b@H�J��b��=����� ������6; ���d� � �5����c��F��4��cy�czJb��f��&��&@y���&��z�&����y&�z&��J��/��� ��ڪ������"=����d��D��D�����"�v���`�����Ϝ�������� �   �i�  5y �v��‖6��"!��h��!���B=����� {�/�����F��8��4��� �&�p ��{�k�(/���@�=������j8�xøK��(��(��&���Dv&,�{���{L�"��"����U���4��b��n\����9ib�{d�~��"F���
.��&��+��!w<)9y������@���i��H �n�l��!��{�/�"��_���A�/�A��|Ź�v�/�%� P�X�c��/�N�B J���|���X� ��#����X� ����1�5A��D.�,  � ���2H����c(��!S�(���N���3��e�/� H �Q��?��"[�"��e�/� H d�/�ôß�.M�^@��; !�@M Â��OH{ �A�k A���AA&��!������?��#��&��Z/ �H��&# ��7Bt&��"�����"���N)$��# � P�Y�cM)$��# � P�Z�nX ������� ���b��J��2��e�/� H YH.
 ���b��J��2��e�/� H �����mr&ns&lq&kp&���
�(� �;5��OL�H1���	E�/�1�����?�C������2���1�1������2���1(�����9�t8	���/�9�X8	���/���1��8�1��8�1���9�Y8	9	Z8	�	����U����1$��>�W8	>	U8	!�	�����/�����/�����/�1�$��>[�8&�>V�8+�D�K����溰O�d�hb�O��[_�fh�����Y�"(��K(/�J��&�ȟ,Z������B�B�-���B���w�b��t��N%��)��B6�|���1��B�����r��bw�n%"��V�!"��[�!��� ��X���dO�����d�0!���&�!.��2�[b!W���U�/�[�D���[�D���� ���G�ڽ F@�� H����@� ������[��⋋e�/�   ���vvbƀލ���$ٕ#����U�k�1�e1)��è��1����"���G1I�Q¨��1���'�2y��?���1���1��<�>1��1��<�@1	�1��<�G1	��˜ѹ5љ��4=��D�b���1 �Ei���6������� ��{����pݧ�� �@i R�H�d�|O X1��
&+���&1����2�6i�1	��(?�:�8��
"ȟ�1@����
"��&Ƨ&1 �1�
�J�D>��&�.��b��&�.�1i�;�?@�1��;C�D(ق������c�M���?��K �(����1���;�<=�1�o�/�;�mn 1��l":1���k:)���<P=<ݹ�J?� ���O1ڜ�&	&�&(?�?�1����y&>y�8�	y6	z6;y�z�	&
&(?�?�8�
y
cz;iyz �"�&+������"

bc���8�<��1��
:91�(��	&��	d�1�����{�����������������I�&�@.HP�������D.��+� � ���ٺ-N�M �F�A�/���A�FKF&��2���1����,�����&�ߚ���� �b		c(��bt�����s�1y���Jy9y����kR�rst�� �{�/���1��9G�� ������ /�{�����{��ﲠ���{��[���2�����2���1+����V�� ��do���O�n`�H�Uq5����hb� �� �� �����6{�/��� � 쀀N���� �ĉt��T�C�D� �  ��qVS!ԃ킕 L� �4�R@ XL ##� p�8vV�C`!�	�� �LC 	Q�TAX��E��GLC U�HRM TR��G��4��AS T ��� p Ň�8�� HR�CkS��H��7VC`�HN�QT�  ��p�8 ă`�`@�� H �R�  XS� T� @��c] NT" �@�g�=8 	� ` R�$= �S� `_ ��E@ҷA- ���T� � �N  T` R�� @τT �  Pσ � ���  �ST�`R��D�MuC��	� @� 0��sLD= ���	q�TAX��E� ���DA��`5� @��tTS	�P 3���T�5(U�AS	�PP@�S�B� Q�u�HRM TR� Hߕt�	5E=8 �S��D  � T�STC@	��R1MXP� P�uC�C� � HL��  R���D ������T���D�` �/ �@ҵT@!�D@  P�8�HTXT@ �KA �E ��C� @�SrɇC �A�4 ��6C R���'S�$�8��C���N�Rנ3R@$   ���B �mH� ����@ �}E���1 ��R� ��	�B@ֽJ� ����@ �}E���� ��E� ��
��A �}E�	�C0�}E�	�B1�}E��A���Π�Π���Š�Ơ����č���������������Ӡ���Š����ҿ�����Р������Ή��ύ����Ġɠ����ұ����Ԡ����ō����Ӡ������؍����Ġ�ۭ���΍���������������ο�����Р������Ή��ύ����Ӡ������׉���Ӭ�����Ġ����׍�