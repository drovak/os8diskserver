����D �B � ��                                                                                                                                   	 	                                                                                                                                                                                                                          �����������r��s���l��� ����Ձ�މ<��/����&�É(Ϩ������ �����Ë���l�<b��k ���'���� �  ��쉜��� �,�볨����ɀ � ���iۀ��!��� ���իM@�dc�T�$���_�9` 8`�O��FE��t?�������ڕ��� �@�����P.�/��K   �&��Ț��C(���������n�,��{ � /������ ���)� ���)� ���)�����'�ɸ��R�t��Cل� @큜�<�r���J��(�޲ށl��<��y����?���&� ��<eP_�T�-VT��P��`��  �
�F����h��R����L�<�b�b��ÉΈ�ww�L(?�ئC���ؖz���������.����L�<��� ���L�<(����h ���   (����6ς �����)� ��d���&��B��   �ز��d� � �� ���É���.����� ��$ゼ8���_�������U��e �   ��̀��  �
���� ���9� (������� ������l�2������ ��l�?���&�'�|���r��k   �cλd����d��6��N�6�B������J����r�����̀3`��R1`6�-T��    ��(����{ ����� ���c�V�4d��B������牬��6��C��b�D����b���� J
�����"��bJ����b�J!���b�?���!���.��b���.��b���Ͼ;��c��&��6��0J��>�ςl��y  8���� c ��L��'8�bH��   ���&���(���cШ/����   8�Oxg��c�Hb��Z�?�t `    	  	                          89I�89I�d
89I 89I	 89I	<89I	 89I	�89I%89I�	89I�	89I� 
89I�	89I��	89I	)89I��	89I� 	89I�89I�89I�89ID89I�89I��	89I�S	89I	889I$89I89I�A	89I�	89I�	89I�I	89I6                                                                                                                                        ��i(����/����x�����r��y���(���c��l��� `����b�b�l�9J
�d�9F�������J   ��s!� ����<� �� ��(��(���@.�/���t������                   6�� � ���U��u���;���`�����f$@���q��n&����� ��b �⺁l��<��/�����B��� � �B��� �l �!��@n��"�����)� ā �� ����V � ����?A q��E3��R���DDN�N	��L@!�O�MN0 	�8��T�5                                    ����Y_ �g ���6�������/� �� �b

�
���(� ���� ��� ���(�(�(�(�/�������� �����o��)��"����.��k��"����,�(/��������*!��&�Ϛ�&� ���b�ӃӝF��/��"�c띓��@��������Ӎ� ������?�!�}] c�� a ��U��Xct�c � �����,c�� �� �0Pr0�) ��9M�@��A%Ѕ�A%Lt@�@	���) 0+N�A�� s -d8K @A� UC�0L ��Kn��Nm@����@�l�T� ��i��bi ��Xp@��u@ee�@ BP����Ư�tl�i ��  H �
��G���b��h�����'�������� �
����i� T�������  �������̀@ � ���d��2����ӊ����P.��/�٨�!���0��O�٨����J�ъ���ǀ�������   ��J�
>

�堮��c��@��b���� /��@� � ? ?`��؇��� ��0 @͏A5 � SE@��D@� 0҅�OB � ��0M 0Ï�C@ � �P � �N �  NB � �S2��0�	5I 0�� � ��0 @ďDA � ��CE 0ҁL�$ � ՒN ����2��@URA@�`NU$R  �N�CA � Q@�`GS � N! @�N��T � X� @օ�OB � ��P�	3� @Џ�TC � �C � ��@ � �	3 P��P �AM�3 � O�0 � L@� ���  �� �NA � X� 0Ł� @ƒ E�!�D 		 � ME  ͒E ���$υAN2 � GS � N�%� @�X� � ��TO  ׀�X�S � DAL �5 � �C@S �� � #��@�P#��@�$ � υ � EO3� @˅�OB � �R@ �P��%�@͌ ��2�DN � �$�� F ��F �� � ��0� 0�	� 0�� @͏	�4 � �A3�  υ� E�A@��OC� Pҏ� � X� 0��� �UP2 � �RE �@MG @�U3P  ��R T�� � N�%� @��F %�� F � �P�	3� 0ŏ� � � Ǐ�G0 � ��0� 0�D  ̏	�4 � ��3G  Ϗ�TC � ��4E 0�� ���LR � X� 0Œ E�!Ɓ� @�� � ��0� 0�� ��DÏ�T0 � D� @�UE %�� @��NB � @V�NT � ��TO  �2���	�4 � �# � ��C � � ��R Ǐ �  P�� 	SA � ண � ;��] � ���� >    � �� `� FR��� L��]���� P��� �  	� ������£�   c �� �� `��� �� T��� /	 � �n����ڸ �����ض��  ���(�� ����.�� ����+趤�  T����� ऍ� ���ʎ ���M 

�� ୍�� ض ཯�
� ྷ�趣��@  T���غ ࿳� �� `    � ��� � ��� �� � �	趤�  T��� �� ����  � �� �7 �  �( 	 0   � � 	���  @�L�8� ����= � ���� � T��� J       �
� �   �"&�+ �04�9 �<A�FK�PU�X\�`e�jn�rw�|��� � �
���������� �   �������ê�̪�ժ�ު����� ���� � 
���$(�+ �-1�69�=A�DI�MQ�V[�_b�gl�qs�   uz�~������ � �����������������Ȼ�ѻ    ��ݻ� �    �� ����������      � $�'+�.3�             DT  �� � PP��@̓0� 48C � P	��	  @B��  5�@P 0� E � ��@��@�DσD� �$ 0��@ � P# A�L	�3  P�TNU$U@��L�	 S��3 �@PF0� @ˋ�ǀ�                  l>�n>Pp> r> t^�vN xN z�|> ~��o� p��o�Po�To�Ro�Vo�Xo�Zo/ � �  ��,���J.
��

�
�ⵚ�ﳠ ��&��� �最'|� ��/�����t������F�⋃��� �� �   � @   �     �M �A+> +�     ��MO�.N   �     � @� @   �M�G��A+>��MO�N�"N�.N%>�   �M�GA+>���N�"N   �@N�@   UTB 8@C�FL�OR�X^�fi�ow�z�̇�̓�̡�̯�̸�����������������������%�+.�8 � �   0�� �   D0RD   5 P@V DP�3         �(���(���(/���H����,�����&������  @@ ?                                                                                                                                                                                                         ��(����@����)��cŁl����d�(?�����b���ŤŠ?�!������>����F.����0��'����(��H�����!.ݨ/���˂ ���ɢ�����]����ɭ�� ����0��(�0�`gEO3� @ ���'��+ c	@��΃����8����P����I d	�� ���b��$@����&��"ȑ���'��"�(/��"F��� �   ���Y������8�G5 E#O�4 �A�s�8�#`EO�4M�T(	#N���3�� R                                                                        DӘ0��]�1��:� �(����bF�����b��&��6�� ؁l��<J
�����b��)��bJ�����)��n�J.P����U����"��b��&��2@������"��càn� ����� ������)����ߢ���1��� �	` �      ��3@           �>BU썈�Ê����
���F`�
��������������������N A�T �B�R@]R0�  ]L  ]Y0 �N@Q�L%@]`GSU �TPBR1 ���R ��3M��ACM�� y� �
�Ԫ�ݪ���� �� �  �� �  �� �  �� ��  � �� �� �  �� �� �  �� �  �� ��              ������0J���&��� � ���{ �	���(����<H���F.��'�������"���믚   �&�&�t�����0��'���   ���/�����⹽�� ��������ĝ�LS!N�MD� �   G���B���Ʒ�}��������� �/�0� ?@���_���8_N�D �	�� � ��/��������  �����  ��� � ��b��r���k ��(O���� ��&� .�/��<�� ⨩�� ����(/�� �� �����ǉ����  �����i����� �  �������  뢨��  ������  �	 �    ��D�G ��2���F?�S3� � ��G��"����Z� �	�����  �	�Ԁ��	�� �� �� ��  (����/�ؾ���(����������  �   ��6��C�b�����2������    ��F���b���k �	�?����{�O�MN0 �3� 0 �               �C^���?�
G~T�����Z  ��������� ���|����� ������7��������&��2����Κ� ��㚣 ��U�� ��ۚ�ӳ�-�����-��� � S	Ut�DAN�!�R���DN(�A3� 0BT��QIu�NB�S�n �LS!ЃE:! �LS!L�TD� �                   �y�c�VG�� ���<�����4���;����P�� ���0�����0��|�>�����0��|���fخ�Κ�������������                                                                                                   ������ӈ>BU�� �����c��/�����l��0��/�������0��'������������~�<������   �� �����                                                                                        ����*����8����y���� �� �� �� �� �� �� �� � �� �� �� �  �� �� �� �� �� �� �� �� �� �� �� �� �� � �� �� �  �� �� �� �� � �� �� �� �� �  �� �� �� �� �� ӯ �� �� �� �� �  �� �� �� �� � �� �� �� �� �� �� ��  � �� �� �� �� �� �� �� �� �� �� �  �� �� �� �� �� �� �� � �� �� �� �� �� �� �� �� �� �� �� �� ��  � �� ˠ �� �� �� �  ۱ �� �� �� �� ��                                                          ��� �BR1   ��h��~����{ ���"��f��i�O� ���"`��/����D.��bH�ǿ��$����"����b�����+         ֽ栐����  ���&��&���&���b��h�b�b��k                                 >H����� �
��� ���6��ǉ����s��y�                                                                                                                                                                  ��o����                                                                                                                                                                                                                                                                                                                                                                                                 �	��?��2�i�������2�����?��������������������?�F>Ȓ���"����?����r(���(/�� ��(��� /�(/�䢠����@��&��������߂z �{ �
�t6G�"�����0�A%ߨ�뮀��U_�[�������#^���"�� ^ ��&ww�{ ������/����bb�b��c�������&���    	�����{�	  ���)���� ��K �(/�񲠼���?���h���h���h�����)�����c��d�<㽚               ���LX�I�<Q�?�$�ܑ��֕ר^�� ff�&�����i�(/�����b�(/��� ��(����/����������"����H.&/���t��������Nđj��� � ��<��������쉜a�܀��쁜 �,�����É���� �	Q � ��������__�_�O���?��E��[��]�$� ��/����/���b�c(��(��Ĩ����>��� /���l��&��9   �
�L�< ���@.�/�F���À+,�������J    !�l�<(���/���J!.ĉ��ɸLs� ٔCX  �O��A3�8LS! �	�������Z� �<?����� �P��DC� �&�)���p.oN�� .�{���c ��&�&t��� ��(/���(����+����(/������ �C��ˁÉ�������&�F���7���(/��� �� /��
�   ���Ͱ�� Ǡ �� �� �� S#����G�ֽ[��W���`�������O��6��)� �����)�������cb�����)�)�)���O� �QN QO�S�8	�d �WTr��8�3D �A� ��`�TB�  �O���4	��`6�TB�S   �6���<(���(/��(���/���É�Ɉ���к��K�A� ��P �"�D��G����������X� ���É� ����'��&��&��r��r��y�������k|����� ���n��� ���� �� /�/��!��&��)����L�<��{ �	���׀��������ـ��Ls� �ң? �P�	�S����5 �A q�TB�  P�	�SB�GO%S P���� ϻ�T����Հ�P�A� X�SO�# ��f�i��/�����)���\ψ����2���&��J�&�&�* �	� ���� ��>�����?�������������(?�ї��C�����0����)�\ω �� �F��� (�޶�؛ ����j�          �<?��U�����I^_W�C���_F � �
����"��c����
�    ���'�� �����B���\����� ��Ɩ��������h�������@���ŉ<� �ƒb�/�J.

�� ��*      ��&����É��(����c(������"����!��?����D�Ǥ� �          �F ��? ��� �������_                                                                                                                                                                                                 ���?�������FN���&��,��|��C����������i�����i��������(���� �    ��� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d��������D��� ���޴ � (����B���ǉ������˛����� ���� 5����� ���ɀ �5���K ��< ���� F�C�A�s �TEB3R �ϋR���DIV�8��4� �A q��@C1	�S                                                         �(�Ӏ��? ��)��7�����'��'��+ ���bg��J� ��]�R1��� 0���R���D�E���PL� �?�4R���D                                                                                                   ��:^���������� � ���� �ᆢ��b�b��ǉ�Ȁ���<(����b��/��������"�������&�����* ������� ���ǉ����/��� ����  ����ӇD���&���ֈ������� ��� ���d�(?ֲ���J �	����$��+ �            � �����`�� GE/�������2�����̨�� 7�����2(����/�����~��x����� ���ɀ ��� �� ���É����������'��'����:��̀`Sr�݀��0�H��A�3�N�G`����d� Љ��Y��A qO�3�T                            ��������%�V]y��� �� �� �  �� �� �� Ѝ �� �� Ӻ �� �� �� �� ͯ Ĥ �� �� �� �� �  Ô �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        