����   B   �� : '> ;? !-?6%&)2?;! 	 *+^   : 
 	
   	  
 *2	,���������                                                                                                                                                                                                                                                                                l @   s @                                          z�HPP   ��0 0 �� T   �I�� 0 DR��` �D;`T` �BC�8LE����@`oS ŒEÃTO�3 �38N�             g  R Œ  �  XT   � ��H�RA  ���K�   � ��HT@  ���F�   � ��HSS#  
�ń�� � ��H��4  ��	� P � ��HN�  T���@ � ��H� 0  ����0 � ��HA  ���N� � ��HT�  ���W�   � ��H��C  ���O�   � ��H� T  ��1��� � �X@   ����0 � �X�E  �  �O�   �  �
��b�bf����i��ρ� ����0��'���(��J�����s����䆂����r��r�bf�w��   b�$@��� &F.� �+   /�i	a>�����Uz|� �TB����>@������y�������B�c��������(����  cȗ���)���(���y�ρ�����(����  c���(����y��ρ�����H����(��  b� r�J
��!�sG�J����������"��������7�?�梕��A|lz ���?�f ������s3Gf����� ���� @�#������#(��tv� ���0��������|�>����>������rd������������� ���l���� ���ɉ ��I� aN$ �P �TUV�C@!�SA�3L����4�SA�3V�L��SA�3���Y@� @ ` u�   �bv�P�Z�o��_1`� ����y�Ɂ�� �à������ �
��'���Z����z��  ࠜ㨥���w��s��r�b g �J�6�&� &� ��?��  & s����=6�/��<�r��r��s���������'��'��'��'��ˏ�B�$ P��r(p�n��s�ge���!��w� � ���{|̀z� v� � �� � �
� �  � � � � � �   � �  � �  � � (     (�"�o��f��f  � ���Ɖ��؁��"!���&������r��r��r��rb=�/��r�|�&� &�' �J�����'���6@ jÁ7D  ��'�_��!�W�f���|�u��V	���z ��&�6	6�6
6 6 	 
 �J����8�(�(�(�*�٘��8ߨ/�F>ȕ��ݠ/�����bgww���(/��(���(/��(���/���������7�����K�'� �G� ������N�/���� -�p�����/�	%��!��k#Y <�����0͎� ��      @ٔ�MA          ��              ����                   �                        ��� S�O�^�UB��� R@� � ����dB� ��(�?��s�@: ��M��hgD�� �����# i�B p�� &W� �?����K� ���i-�&��C��d�h?��@��~J.

,��2�8b�}id @   ��΃ ��⪥� %�%�&�kL#� �G2N  �R1M��DR	ϋ��� 0��;��R��C ���!�⠺�����ھ��F.������r��/��朂� bx�/�|��خ wb�n��u(����}�ѶU ���ƀ�6� N��6��F ���J��:��N��c

�
|�(��{| {�(�Ѩ �    ���������6z�� �0b!�i�>�;<"F�����������C         &!�̀�� ���(��(� ��zɁ]�yٴ�MA��� 0 X�  �ES3  � b����naih ��� ��3K �� ��l��&Ό,��b����ۊ��6���x(wߖ倄���F�x� �cրd��6��C a.މL�0?���� �`����㨺� �� ��� � bJ
�
��� n�d������؀c �'������/yݹ    �
� @� �      �v��  �����&��6ݠ/�����b���� w	��&������}?� """Bu�~""ts�" & x0 ��$�k ;�ͨ������6"  bc  70�"0�j�Ǌ0r �0&�/�~�66&����q)~0"~p'&@>uo %�&sr&����/���� ���C(��<<b!;��/�͔� ���&�<6<!.;�b�g��{ �
 X"'ӛ�t�O\�'e�'�hgD}�G(�* A   � �

�
|��&(?���n b""ca㠰�"D�J�"Cx$�"�t"�

���'cx!"n0"�{���:7' "&��"7"D��&Dn"��/�v��� "�"�#�k n&�"����?��K >>�9>>4|��m�m�����7W)V��7 /W\�(7���@U�Y ?� ��(?�}���<�G ���x���r�b!�'�(&�+&�,��=&�2&m������(�b ��(+D�����+b(����>.b��(/�)��)��)�)2}"��������c��G w	������ �b

�
���(� �| {| {)��vƐ�*q��3��  OT�08D�B7 N� �aFA ,� ��=�=�n,�h==t�=�=2D����=&�2&� � . � o =�; �}a�� � �� ��>b�b���bn��)�J��� 	��	�9�J	!6	�8�!��� �l �<�!����{)事   �>�!.��>!b��׋ ���� n ��)>&	�8ꀰ�� 0����
cY��0�i1!.(��1b�hs"1d����������&�7�7�|����c��B w	�������y�����; @�󢱯j�vy5�Q P� @��"�i�"�q ��$���''Á�"o F���~2b�|8�0]Y�\�"�"։lց<$���;� ffieF � A1�fd�OR[�$ ����q)#D 6C b3b4�h�bq-�D6&l���?���k�k؞74�  bo .��#k��&2tk9�� �6t)#a>&� n"a> H/�H�.�b##C9#d!.#H?�:����85�kv��ó�$t	c%� �)����ɥ����5 �8  m	��)�	&	H?�!�{)�!��m�� ��&��l} ��  �� �-.  c������-(?�-��v�-�P N E� ���� @�)��*�@&�*&%�)n  )bj k�k�� �	  bu''�"cii .�x���k��� ���g{�������j �)|������ a����;�Y$ -c!9⨴�-�&--6-.��c!9⨯�-�?�P��?�خ�@�9�'�:B�~��b`9␬�9�&��/�-� ~-'��� s-�&��08�c��Ѷk    �/�7����7>X7�� �5'�5�8!.5� ���9~"9:b:&�8�5�k P��/�󩀀�H����H��7��H+�E�s�8���� �	�̪��x � ⠙�ဎဎ�k)�k)>X��� �/���0r cr(�!� /�0��!�/����%�jj H4��~3�'�h)�)�n(*�/������'�/���'!.'�hk'�ρ��I�0!0��(��7f� �2�J�}�   �+&�2&�+É+�� �ɔb��G9jTk�@��� Ne� �q��� &$�"H��~H. �0!����l�<�Jn�� `���� g��f��f��f
�;�<�&�0�, d�0 '���ti%�'�y� �ki���Neimi�ki�mi�mi�m)�Ei� ���?���� ��"��Л"�(�U�8C �R1҃@�R	A�1�8I�PH�� + PU	����!�n$(/ݞ����r0! �0r (�� �/���!�$�"  k���ݣ�����ڪ�0�r��g� fc@n#2f~" 2g r"r#r'�p'&0�*0r ���'h9�'� �n (?������@&�##7%�n""�z�J�JB'��'&$!"iy 'c��" @O頮 F."�%#s&�{�gD�~���kG�t���������Ψ/��b�i����&��f+(f�	��	�i�J�/�Ш"�n �l	�< (���?� �������c(r�s+'1B��i0�is"�b�d��� 
 ����}�z� ��!.� &� $����&��&���	�l� �      ���
�|z�e�r ��&[R�/���q~�tBF���li��H>������.r�/r�/r@u�o./F�2���'�&���'�.�H/�� �� ' 2"2�e��$qך��!> cnF�72'5'5 $һ� �&l��i%�j(�"�"J.x"��t)#@>&&7%�n"%�zi�2!�X(@�*�0;)� #�.�'/�',(/�0����<�lvߖ�q)��v� /&�����|C�t�7 �'���}2�FX������<�B �2�P�⸼�v�2�'�&��<x2'�'�}�d�H� ����	�bjb c66bJ�n	6o 	s	s	t �J�6&��� �      ���c�&kCA����6V32�F��� ����/��������j&��� �j�&&l���#���i&��� &�y."��v�   i&�oD%>5�&@>/>&/&'>/&%�.>&>j ���.%'>.&� �g02fsgrtp�h՘#"w� �"a>%�?�#�a&���"%7#&7� ��	É(�� �(+"+ b(�k l	��xJ���� )�����L�����{# P��,��l��0(��J��F.����& � �术'8� ��/�����t����  ��� 0�ob b��bvi�#�b#%6�!.#(?���%!>��/�%���J�v)T�&#!>��?������ᠮ# 0����#�##s�%&�%'�!.%�"�S���b��f��&C &~�*� w�q��? �O���Ơ������Рɉ�����ӱ������ō��������֭������Š���Š��Ҡ������ˠ�Ơ���Š�΍�����٠��Ġ�Ϡ��٠��Į����������̉��Ӡ������֍������Ơڱ��ڱ����͠��č�������ұ�����Ҡ�Ơ���Ԡ��í���������Ơڲ��ڲ��Ϡ J��J
���
�l
�<��|
�<��s����É��J
���#��� ��J

���'��0F��⊞�JN�FB�MR�A�MY�JN�JL�AG�SP�O԰NֳDC��Ҡ����Š���Š�Π�����ҍ����ĉ������͍������ɉ������ω�����Š�� ? A@K�F���dP�@�?�M�