����   � � 4	83
4 ?2?>4>?<  =9	2=425.=?=>=7=82=.)

:   ?=0 =2=3=/> == :���������                                                                                                                                                                                                                                                                                               �h��       X                                  ,~�/%˃}�Z P       �  ���`.�Q�� ���� �� '� � �� �� ���R�q�^ "
����x�"� ���t� yrt/�n�~w�x��n��" �p �rs�o��}�� |�{c�b`z���d���zr{�~�+2�j �zyr� �|!>xx7x(?���!�n�	�w
&	
7	"����z�y{'� ����v	&���v
&�	� �l
6!. �/� � ������	 6 " u���" u��� !.�/� � ��/��  ��/��K �f�tɉt��K��K |!x㠨���	�n		r%h	�Hs�"�?��		r@r␠��q�R���xTp7�Lo&|�[ nme�l�����k�l�k�v�j�m�in'�h�� ng͚�f�leUedRgmsDm�} m�zgH?gwc0Dg��@n�gsb a /` /(�_�(��^(/�]� \��kp�Zl�^m�{[��ZbYX�Ӂ�W��W��$�VɉVɁ|ǉ|�X��U��$Xi���||uUژ�|�!��|�?����|�|!>�|è��Uژ�|Ŭ�(��Ёl|�<�|����!.T�& |�`x㐛�|UY�Ɗ W鎁�|�<|�?SR� �|Q7�|�Qr�jX�U��ڋ�J�S�PO)� ������ |Qc|rQ�{ NM���L�҉��N�M�� |!�#�lJ�KM)JM).�		cb!⨹��&&�� �j d/@����� I"M������HM)#G ���	(?�m�(��FM)�\�MN�M���� EM)�J\M)NM)�k$�J�D�Y��CbMB�M�胬�Ѱ�/����J��q� 	��&��� � A "#d�o²�l
.���".c�!!7"
.
�c � �! d" '�J�Ɉ � �
����@�?�ZV�q��� >=b �k <�/�/�;��/���?�	���c: /u�/� �		& ��z 9 >S<�n98 >7:8c6�8�5c!(������ �� �� �� �� �   	� �@ٔ�MA��;�!� � �"                ����   �L� �   �� �� �� �� �� �� ��    &~>&}&�>D>��|Z&�Á(�{��z� ��y xZ.
�Cw�v'Nu'7K ���� �� �����6���2��}�y���� �m��/�Lt��/���z� srbN�l7q�N�l7p���lo�< ����lz
�T � �
��,o�z�z�  �n�obmb��l?�D�٢�b(l�oc���z�   芬z	�ڋl�k'��+ي,t��oÁz�  �
�Lj�<�i�� ��J�n�hg"7fb�7��e��d��7�����t��
 &!�ʀ��