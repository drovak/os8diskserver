����  @>?.8'7/'7.-      :   :   :   : ????????q7,<,.).  (/ A3������������������������������������������������������������������������                     C	D@�������%!.cq9|&R!q�|o[� �%�&-bp(�b)�w$��
(᠐�(�?������)k F��!.(/�!�&���a4>X��8+�`&����?࠮&_&&$'&'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?����`!��k�\��l)�� 0[�   �� �� ��i� �;`.            H �                                                    � UUU(/U6 W71wI�w� V ���p^ x  B ��@    
/8��A�.���������]��?��A����2�  ��������/�%`�,D򂜪YɬC	�b�ZV���b�b��b ��D�C��b�ZV��5C�bZ����  U
U$+U2�WAN2�8D��!B � (/�x�(w�v(/�u�(��t�/s��r��q�q'�!�s��&sK�*!��"��*p'+o',�+ ���f�h���n �bD�.Hs�b �J��"�*n &��,�/l8�9��/�����?�r��@���/��8�b���?��x��@���/��9�b���?��x��@��/�n< �;��/�?��x��@�����7� ��/�?��x��@����H� b����t����s�c�*���/�-��b�p�   �
�@.b/�F�u��#��r���"��/l.f�&�<���6�:)b!⨘�?��~��A����J@��/l n.�b�b<��6)b:�!.�/�?�
~��A���D�J@���/���&��%Di��7��0�/�?����A���D�@����0�/�?�!������bQF�u�7� �P(/i �Oy��m�L# /�/Rb,�b+�bf,�<��=V�Q2;)8�!.�/�?�;���A���D�@����/�b,�b+�bf,�<��=V�Q2;)8�!.�/�?�F���A���D�@��̪/�b,�b+�bf,�<��=V�Q2;)8�!.�/�?�Q���A���D�@����b6�ʀ���������/�b,�b+f,�<��=V�Q2� ;���;8�b!⨠�?\����A����@����/,f�b+�b�bf,<)�=�VQ�2b;�;9�8ib!���!.�/�?�g���A���D���J@���߸�(� �e(�>�e>�ߋ ���������=�(�(�u� !� ?�?���/�b,l�b+b)&fVP�33b���/f�/��1�E��&&,<)=V�Q2� ;���;8�b!⨲�?-�~��2�/�V�R�_A��V�O�����J@��12f�!��!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E �?��H��2�1�/�C��C����1=i�<)��+&� ;8�f����J+&.�;	���V�R�_�� >	8�E&�d��� �Ji�!�V&r�B��>�bWr�c�t�ʫM�� ��ݢ�!|�ԫ�����d��6� � � �ۢ�݂��d͊���  �������J� ��w)  J
�
��(���2�?� /�b,l�+&�b�n�&b)b*'f&ViP33�/��/f�/��1�G��'&&&,<)=V�Q2;);)9�8 �!.�/��! ���?4����2�/�V�R�_A��V�O����D���J@��21f�ز��w�b�$�8�� �8�0�P/A��!@��������}R��_�=�O�@��2�1�/�C��C����1=i�<)��+&;)8!�9 �����J+&;)���V�R�_�� a	 >�8!�9 �G'�&bd��� a	 ��Ji���}@���lt�$$bp ��X.��/!�x!����"k0�!'$�J'j;P"F�i�h�+Ii(g�**bf"&*e"!*bd(&!�;�ӛ����;��<�T��B�@ a	 H쀀�� �a �J�_�� a	 I�_�� �a �K�_�� a	 -�2�/�-�L�˜�K a	 M�_�� �a �N�_�� a	 O�_��,�P<)�+�-bL �4>i�J�'�'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[�   ��  a	 %擠��%��.�����/%A/��� �a ��%�(��DQ��Q��AH��`�00b5�+ T�$^)�&�v�,.$T�!_bU`�!�S�/R!��~!!&��!bq*⠽�_!&*&$^)$t!�JQ7U�rP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!!.��� a	 ���&H&�&�&&/A���t�)�J��F?�&H.�b'f�A�D>?�'�'d�A�''&&H.�'&)bH)�O�3���������ŉ������à�Ϯ��������͠���ō����������������������������������������������������������� ���� ��&'� ���F'r����'&� ����)rJ��F?(�nA��D����((&�A��D>�/�(�(AoDP���((&&H.�(� A&�'.H���(� A'�*H.*)bH��� )d��3�/���_� � ����Ԡ����Ġ����������������������������Ġ��  @  � ���&V�������6��C��d�6�/B��� /�B)C+�C �C �J����"�ViK����_��� �� x  �   VM����� �VN�����V�S��C�EUy����'   %%b��%bӮ�� ��AF���A����+ ICi�sBC�,t�ޫ������������í��Ե��0��?   ��6�CA���A��� ��(���H����* ����� ����*�^)���� p������͠������������Ω���������������������������������������������������������������������������������É������ïظ�����������ފ �� �?�          B    BĠ������Ω����������É���������­É������������������̠���ԍ�������É�����������É��Ÿ��а�����Š������Ҡ���ԍ����������������ŭ��а���а�����Š������Ҡ���ԍ���������Ã� ��A� 5�A� A�	� 5C�8R0D`�d� @C�8R0D`�d� @C�8R0D`�d� ��t OR �P	��4 �S�ϔNE%� p��t �P q\҃R�Tl&=V�N }��,��D΃	�S_���t �T҃N� �S�ϔNE%� pC�8R0D`�d P��PR��H�= �@ �U�R��D�} ĉ ��PR��H��S�D ��PR��HRT �� rȒ�C � �v��� 0�� ��� SD��C � ��� D0��� 0��  �� SD��C � �rT��� R��D�� v�T(� 1R���G�5G� �'C� ��G2 Ʉ` 8C ��pR��C �NP�TB Q�UC5  ��@VD! �NP��D��NP�TB Q��@VD! �ɇC8CcÀ1����D�4��sG (�FB �T` 8C ��t�3C�8�1����C��G�G2NL   ��FB �TU3 Q ���VD �W> nb����8� D �����������������(���)��������� ���/��� �榤D�����K      �m� �D  ���� �Ȍ��+ ������s� ������d��0(��@�
�

��ܓ�(��@����)��J   ���� ���&��'݇�@R���D�8TT��@�?����� �����  ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    �
�}�to�nm�{|� �����Ъ� ���r��������i�����g��π�ܠ/����&��I������   � >��y����������������������8�e���@����»RS� Q̍�������6��H��h� �   ��)��9��� ��?�>��� �������)����������TN"�  �	���/���g��)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP����û ��8�A �QS�R���Ļހ
��i��� �F��b��b��Ė�d���    ���(� .��bĥ����   ���A����������� ��� �	�Ô��Æ¸+    �֠/�բ&!��"��բ��ز��� �   ���ձm����J��J��6��i똸�כ  RQ��DA���8 �RS�Q���� ��� �� ��� �����A�����Ѐh�����������:��D�����G�����J�����M������ȟ������ȇ���'�Л����m� ��C AT  �� �C� Q�� 茀���������@	DA�0��0,�� � @` �� 5N���@1�N�� 5�N ��;��A�� �/ �I�3@N���Ca QN%�PE �SՅ-ORQ��5` N���N N�TP U��0� A�Q`RQ�4N %�T � RC �TNB U� @����DN"%S� �T�0"��CS���D�0O�#�TBȠN(�U�$5�`%6 ��RB 4N %ER��T �C`�T �