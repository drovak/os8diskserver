����  � 	  		 		   ;   8
8
8
"+ "+ *"  ?<(.	>>(=<	#.+  : ;#:#.8  : 9#.?  0&0!+: /  00+0/
U9 
     ?6-���������                                                                                                                                                                                                                    �@ٔ�MA�� ���      ��� ���   @i �  �&���(ˁ��d�� ��8@��7��@� ���Ѝ���"��"��"��"JU8?UDP            ��              �    �����s�
��� �v���? ���?���R��` ���!��&���&��ff~$&ǝ����������i������z�@y␪�x"Pw� �Ed�d� ���d� ����e� ���Z�Z�"���Ƿ�Z�"���� �������K �b�k �BO�F֞Bc�A��OF)cA��b��
�

������ u (��|u |)�ظ�|�3}/����  � # �� TTb!S����T�S�n� MN&N�0�U��N���R�n� 
�RR&����O�n� �a��a����U"P�n�/�U��U����O��b����a⨀􀅴�e;SWn �� E�pJus �խHt�c�%\�� �AP�Cr�   � `� �  �BQ�DO�PF)RC)cA���� �OP"FR�Cc�A[��O�P� F��Cc�A[������K������̀@ �����d��2����ӊ����P.��/�٨�!���0��O�٨����J�ъ���ǀ������D� ���J�
>

�堮��c��@��b���� /��@�v��?�?`��؇����� �JH�m�(��� �WV&.[�[Y XL)[.[�V�JKK�� ��W�V[fIZ��Z�Y[�[Vd�[�
�b�H�pJ)����_��Z�LZ���/�Z���/�Z���/�Z���/�Z���/�Z���/���_.���Hr�J��Ht�J��Hv�J���V���/����Ҥ= �� p� p� p��HPs�nk�}�����������b\�b]\c^^c�^\t]�JJH���)J�����"��"��"��"	�V�C`!���@N�   � �� ��ڷ ��� �� ���� �� ���� ����) &�)�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2���� � JJ�H��JH��J9JH��J9JH��J9HٓJH��J9H�JH�.JIHL�JH�dJIHu�JH��JIH��JH��JIH��JH��JIH۔JJ�H��JJ���D������>�*�!&�!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0��0  �  �  �  �  ��	��  �  �  �V�3��    �  �  �  �  � ��5 �LG�N1 X��AM  � EPX�U �$��R��A�3� @  �  ��0r� =� ���E# �0w�@ �  � �� 3X  �= �0-�	���5C�  �  �  �  �  � 1�-��LB	5�8E��E���d�����    �  �� 4 � =� 0�-�LC SŠTD ҃	��E� 0  �  �  �  �  � 1�-�LC PU�DD ҃	��E� 0  �  ��9q�`=� ���@���KA/�	�1��  �  �  �  �  � 0�-�L0h    �  �  �  �  �1-�  �2 �  �  �  �  �  � 2�- � 4�    �  �  �  �  �3-�  �v �  �  �  �  �  � 4�- � ��    �  �  �  �  �5-� 1�5 �  �  �  �  �  � 6�- �22�    �  �  �  �  �7-���L�N!�OF`Q�D NRXà;� ���A��C`	G��CBS�`S#L�S�8TO�# N2��TO� 0���`�d`
>

�`��`�� ��(�\�\� ����\"ī� ���(��(� ����Ŀ� &!�ʀ�� ����l�&��&̥&@��tO��t���( L"�|���� ���g{�������j �)|������ � �� �@  ?                                                                                                                                                                                                 