����   � � �� ��>
5 ?     );*A?+2$��������������������������������������������������������������������������������                                                              ���ڰ������������������������������������ڰ������������������������������������ڰ������������������������������������ڰ������������������������������������ڰ������������������������������������8�  ���  0֭A�	��@�EE��� P   �� � Ʈ "4="��!!� F ֔A��PP֔A�����֔A���� 0֔A���σD֔A���P 0֔A�B��A�|A��T�DK��� R֔A���  ֔A��� @��E�����ME�C�	 D�J���S�TN*���S�T� �@�  �� ��������������I���)�����!���K ����� .��d��J��d� �    C �� H �" ��/�� ������&�+ ���6��C�(�@��

�
���0(���@/��"�� �   ����� ���&��'�ӳ� ��
�����@�?�� �  � �����;��A����b��c(���/�����J�/��~����K�B��}&��"��c��k    3<}tq�on�m{�| �DgmJNYr���w������f����i��w��w��ˀ��������d����� � � ��������� >��{��y����� ����[�"��"��������6�I��h� �   �))� ����������; �� ������������TN"�  �� ����/���)�)I���b�i��F�&��J� �!�����"����"���� �k�)��疮 � �` �� ���� ��HP��� �R���"�  F����&�� �)�.�撆J� �   ����� ���)��J��   �|�A�|�������� ����� 	I��b� �ځl��<��c٠�۲٠�ڢ&!��"��ڢ��ر�ڲ�޽ �    "	 ��    � � J�~���#�;�~� �	ӄ��{
� ��"ۊ �� � �l�Ao��n��&� �����?��ƒΒ�)ђ�)Ԓ�)ג�)��ȟ�!����ȟ�����y����� ����r�r��s��b���   C �LD  �� �C� Q�� 茀������ ���Ȉ ����   �� �         ��! ���   � �;�,                                       �
�������������������Ȫ̀���͈� �`S��kX�1g�!E� ���Ι׏���  ����������������������     ���݄܀�̂��    ?   @ �   $ ������ �  S�������3��5��b��L�5e��b��F�`�5�����M��5������N�i5,�����O��&&O&'D���5I����5B�����]5S��b��(��!�(������ i��m�i�j�i&5]��b�!!b�/�!��/7��j�����'lkf��/�s�\�)��8:���0�:�� �Oa	 �^�_.it-)��8y�:���#��8m�:���%��8m�:���&��8m�:���+��8m�:���,��8m�:����0Ґb���9r����:����/Ґb~�/�9�r޻�:���� ��2���� ��W7eX'G]�f]rgFy(ؔ� ����TarU'y��Kb/�F�u��#��r���"� ��o&fy&b.0�/ib!⠗��/�9�r��>����p"bt&�J:���$�.0�/ib���~"���9r����:���fybf.)0�/�~"���!.�/�9�r��>��Īp"bq&�J:���$�.0�/ib���~"���9r����:��m�L#� � N�{o"vb-0�/ib���!.�/�9�r��:��$�0�/��/��~�/�9�r��:��<�o��bsb-;�;0�/ib!���!.�/�9�r��:��$�0�/��/��~�/�9�r��:���� �`"��b�b	�b `F9	t� ���{���������A&(?�6���$�v-)��8y�:��{-)��+���+��8��:����8���8����+��8m�:��v�-$�+��8m�:��$�{-)+ �iH.�����,Ě�,��8��:��ʪ8���8�����i����$t�-��,��ڪ,��8��:���8��ں8���,��8�m:���� �Z&�2��J����(�u� !��&��<�� n<�?��fsr-;�;0�bu��9�r��:��}�-;�|&o&0�/�!.�/��!⨰�9r����:���W�b���9�� ��:���f�Xcb!���9�����:����&ؚ�&��8��:��ު8���8��պ�*�Xcb!���9�����:��&�8m�:����@���E��� 0� >=W����8��:��<?��|�-;�;0�bu��9�r��:����-=�=W����8��:���^f_Lb �f[ .<i?��G�fFyZ&^b.��}-);;�;/�o�\/H.A��J!.�/�9��3��>�ᳪD����^q"^d�J:���.�^_fj�/�� �Jp�������(��H�� �<?��]�f}r-@��0�bs��9����:��)�0�s ���9ě���:���[ .<i?��!.]�/�]���f�z�f�g'}-)@��0�s ���9ě��>К���J:���[ .<i?��!.]�/��g}r-@��0�b}��9����>��ժD�:����              <?��}�-@��0�b}!}�/�9����:��)�0�} ���9ě���:���[ .<i?��h'}-)@��0�} !}⨼�9ě��>Ě���J:��� �                                                                                      <?��}�-@��-��'�0�v ���9r����:��<B�C?��A��}�-@��T�b���9�� ��:��U6b&!.�/�9�����:����%��Ī%ʚ8��:���8��ĺ8��:Ě�]�bcb!���9ʛ���:��0�� !}���9r����:��%�8m�:�� ���D��D��D$�؅� B<�?�� h�A��}-)@��T6�/�9�� ��:���f^_fL .Ci[b �<?��A���hHybcwF��_.)�}�-@��H�c6F�!���9ʛ3��>̚���Jڠ��_�t_&D�:����.^�_�j�S0_Q UX GM %��ť��U�oUm�5��U��U��U��U��U��U��U��U��UY >�[ .CiBr�!�gbbt�<�?�A��}-)@�D���9�����>����D�:���� �]"(��! �PQURSUPQURSU���]�/������ ��P�QRwS�{�������͠���ō�����������������������������������������������������������������[ .CiBr�!�gbbt�� .[�J<?�A��}�-@�D����9ʛ���>�����J:��K¨E�K!.Kb!n�O&[ .fC<�?��A��h'v"}r-�!]���WTU@���@��-�T >���9Л��>����JD�:���������������Ġ�����٠��� �K�!�K!.nO"[b �[b �Ci<?��A���!⨵�!.]�/��hrv'}-)@��-T����9Л��>�����JD���J:��<C�?��A��h}r-@����#��Ԫ#ך8��:���8��Ժ8���#��8�m:�������ٍ����������������í��Ե��������� �K�!�K!.nO"[b �Ci<?��A���h�y'}-)]!.�/�W�T@Y���@��2�#��9����>����D���J:��K�!�K!.nO"f[ .f[ .fC<�?��A����!���!.]�/��hr}r-@��2�#i�9��&��>��̪D���JD�:��E�����*� ��6�fBab	c	cb!⠕��J���� �Z�;i�J�.� �� �a& e�	sb!�	w�J� ����;i;;�=���������������É��Ÿ��а�����Š������Ҡ���ԍ����������������ŭ��а���а�����Š������Ҡ���ԍ���������� ��6�C!!b��!�(� �m(�z�H����* ��� ����*�4)����� �  ��㲧d�"6��N3i xabg�J"&a&6����!�"���!4)!'D�ᩯ���&(?�!�����J�6�������� �
`!� ��!�I�!�+ I	��&�!���������É��� �@7��H/7�� �a&!.f�8$��F� �b˙ �Ϫ&y&M"&��� " �"D��� �Ъ&y&N"&��� �"�7��"�7�� �H� ��-� ���فz�������������������ɪ� �55��b�K��¹��˸Š���ˠ��������Ҡ������͍���� �b6�#�7��"H7�b�!.Zb!(��(����7r�qm"[[b H�[\��J ����4����&�ܰ ��4)��� �3���޷ I	��J�q��3�����q    � �^
.�� `� ��_�

�
�� `� ���� �c��tlkf��������Ġ���Š�������ҍ�"�G	 �� &��6��C��d�6� Nl�h k� ����Ju����k�/� ��3�W3� l���3 �l�/�̨�Jiv�� �I!���� �""b���"b�چ� �mAF���A����+ �3i���3�X��̫� x  � �0� J	t��k��II" �� �k�/�J�r��k���Js����� �������  �� ���� �� �ߏ�K �� ���� �� ���� ��� �	߭�K 
���� ���� �� ���� ��� ����s���� �`"��c�c	�bFi 0	t���`�"� `��񀿂������'���������̵�st"�q-A�Š�	G��4C  ��tC�@޷���`1S �O %�-E ����`1� �O %�-E �C� �H��@K��pRC �T��@�TO�# �كCăm ��pRC �T�3@[��p�EB�G@�O@ޕq8PS- `�sDRE�@;�GT� �TS��� 0N%�PE CP	�U �	��R� K�PB N�TP,U���PB �	��R� K�8� $τTՃ�8�08 � �NA DPS��C �P�CA UN�R�DS�R���D�8��C X��C �� DR��A�P��� 0 ���D ���D �S� S�� H��D ��� @ޓt� H��D �X  ���� � ��� @�q XDP � ȀR DP � �  XDP � ȀR   �D  �Xq  H��@ ��L �������������������������������������������������������������������É������ïظ����������Ġ�������� �������������������Ġ������Ω����������É���������­É������������������̠���ԍ�������É�����������É��Ÿ��а�����Š������Ҡ���ԍ����������������ŭ��а���а�����Š������Ҡ���ԍ���������É�����������É��Ӹ�Š���Š������Ҡ���ԍ��������������������͸�Ơ���Ġ�����Ҡ���ԍ��������������������Ǹ�Š��������٠���ԍ�������É�����������É��и�Š�����������Ӡ����͠���ԍ�������É������ ���É��˸Š�������Ӡ������̠���ԍ�������Ɖ���������­Ɖ��˸Š����Š������̠���ԍ�������Ɖ���������íƉ��˸Š��������������٠������͍����������������ĭ��˸Š���ˠ��������Ҡ������͍���� ��D�J
�
z෧h�C������&D�&FG�@���F�D�$� ��L�D�hA���L����� �C��@���o�D�DD�D��D�d� ��A�񷇁G�@E��F��D�� ���K��"��k��A�Էb�E��F�(�!��H�zJ��N�����N񘷁<�Ř���E�   ��       ��U�0�H�� I	�����I�����`v�v� ���c��d� �����+��L�'�'�'�'!� r�'��'��,� � ������'����{ ��<  �    ������hyJ
���h�F����i����,�|FG�@E�� ���@�D�+ ��h	 �����7��� ����    {�����