����  �*?9  h<> <(''%	$(	%)( ' )				"#						 	!	"(  /'<=';
:<<;<8!;> <;<'+//$    )>B   j 8? *
34
5
6	
 	*��Š�э������̽������Ơ����Ҡ���̯������Ԡ������Ġ�Π�������ō������Ľ����������Ԡ����Ġ���Ġ��Ǡ�����Ҡ����ˠ������ũ�������ӽ���������Ҡ�Ơ����Ӡ�Π�����͍���������Π���ˠ������Ӡ�������Ġ�� �C� � ;`.  � ���/   OQ'PR'��pl5'�/H�Ib	6hJ&K	&6�MN�4���4k�.� LSc	St96�����;Pܺ���P�=�B����������  ���`��/J�"�
�F��! �?��A����2�  ��������/�%`�,D�� �(����'��J   � ��&��&��"��c��s!��� �� n��&��J��    �������0����0�����7�������������!��?�(���7��/��� ����Ԡ���b���&� � ���������6���� �hd'6_t�a�fg"�&hce~* ����!������s�����/����!.��;�(ύâ�����j�����/��"��l��"��lֳ&��&��6��6�?��s!�Ġ?����J��B�o��  ��� �������~��s���� `� �� ���c��&����b���@���׫��ɂN�e��U���"��"Ā �� �dԥ  �����"H��q�☈������b�&����r��n�/���&���~��&�����~��(��'�D.�/����&�/��������b�&����'�����j ������b��r��r��{�����)��9��)��9��)��9��               �����    ������%�JTW�D ���� �� ��s!��H�����(����b!����y����y���~��y����y�� ��)�����0��i�Ś�Ś��|��'��0��������ʚ�ʚ�ʚ����/�����/���H�����끼 8	� � � � � �         邐m�S�hi33;3H1�������� ����1!�����!>�?��!����������!>��?����������!������7�!������7�!���?������!>��?�����y!���:���!�� �������ɂ�����������ʠ��3� �逞�(��>�e>�艂	�D;eJD����Q���fg"WU��� � �����F.��b
����b�����9��9��9��0�����7��7� ���b�@.�/���!.�/�q��/������� ���c��h��B� ���c��h��B� ����!��H��q��������� �D��b���� J
���&�'Ҝ����     �    8������e�A�d���  � ����'����'���&��(����/����s���0����;� �  ��  �����'�0����0��/�ƪ�0����0 ���죭���7��7��7�����|��'�0����0��������8��8� ����ኼ炐D���Q���fg"������U�D��A��U� P�򣹠��s����s���򓵠�򓱠�򓲠�򣴺(����/����0(���(/��������2�o��   @ ���� �����s!�����!>�?� ���&���l��&��� ��?����� ���'��� �"�i�Cc{*��D�U��U"1U?PU_�U�Q� 㩦�0���扚�壤��穐���0���藚��C��������0����@�  ��   �0(���(/�Ų(���(/�Ų(���(/�Ų(��Ĩ/�������9��9��9��9��9��9��9��9��9��9��9��9��9�� �	����U��U�,T��U��U��U��Q��5��Q������Q� 0� ���&��cD������$���D�杆*��{� � ������{  ���Z��� ��>��&�>��J�~��{� �������c
������ ����
�
����������� ��>ޕ&�>��J�~��{� �������c������������/���������9�h��� P� ���㓓d���� ���0��&��J���� �� � �����d�����K��7��{� >����{��6��7��'��������{��7�����w� ��n�l��o�o�!>�/��!�����!.�/��!�����!.�/��������� �          �  �1�����6�t��U�,T��1�  �����c����!.��s��������'��)��� ���y�&��� � ������������'��]��¨/��C�����U����'��'��&��� � �����6����o!�������_��B������D���� �    ���d詂,�c�R�6��f��f����fe� �W~���, ���������"�à����D�����b��i�&,���    � �^l �㨭�]����� �CB�A�������/�������栗漻&� ������ ��������b��d�ڤ���� ��?�>���� � ����b	�l��&�Á	���J��� �k��y�	���A�`�b�Y&TU�S �� �����������������I��&�/���)�������� ���/��� �欪D�����K      
X� �� H ���?��� �������'��; ���6��C�(�@��

�
����0(���@/��"��� �  � �?��@p�+�$��=A�	���`/6w�F����ƈ� �� ���s��������A��v�&�(?��������D��������9��)񁔁����;��2��r��&��6� �   }t�qo�nm�{|�  �@ ��g�ϛΠ/����&��I������   � >��y������ �������&� ��!�傐��w�Ї־wX�xƔ�.=w�SyUT��ň���ghb p쎨��/�����d����    ������  � PH�� � ���㕨��i��������� ��0����/���&�i���9��)��Y����r��i��F���7��J� �!������2�����2�����0��{��)����疬 � �` �킐�i�.�p,ƈF=w��x�����x�\i� �� �Fb��b�����d���    ���)� .��b������  �� �  ���A������0������� ���I� ��Ŕ����ŖĻ+    �ڠ/�٢&!��"��٢��ر�ڲ��� �   � �������TR	�S  �             �	����.�x=�w�S�UT�� `� �����A�������cר�������钖�i>꒚�iFҒ�뒠�iIӒ�쒦�iLԒ�풬�iOՒ���ȟ���ȁ���'�қ�
X� �LD  �� �C� Q�� 茀������ ������y��{F�HL�NG�I����i�>	FI�LO��F��6�І.x��x�g�bg  �� � ���������h��J�����   &!̑"����V0���++�D��,�(��&0�!1�0j�+�(d' ����+�� �@�����P.�/��K���b�nl0D ���2� ��'D���ᠮ# 0����#�##s�%&�%'�!.%�"�S���b��o �0�
F���W� �`������b��g��6� ���t��6�����D�Ч��y����������{��#��s!��H�����!��!�Ҩ?�ҳ�����7Ҩ?������ Р?�(/��&Â�Bf��`WdBhe2W�h
�@�� V*WX"YZ"��3[\"]^"_`"ab" �����&��&Ӻ"��c��s!�����D��J� � ~0�.�����'�&�	&�S&	7S�J��'���b	�bSc	St���
�����J��J�Ι�f���� ��@������j�  ��K��&����@�����º��P�E.&F/&D&����D��i7�J.8&/9&8.&9/&CCB��/��(/�����z��j��(\T/���� ����-#�%� D� �/