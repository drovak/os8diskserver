����  �	  	   	? 0= 		   		    	     ? 0=     	                                                                                                                                                                                                       ���i �9"`8�    +��/           P���� 7 �� ����r	  @��b("�jb5a��� �  ���?��!���Њ� ���@� ߂ 4!Ҫ� #��W���`� �/K�"�
�F���� ����V����2�  �����"�/�%[�D��D��D����9��9D�i��9�/�����9�/�����7�v���l���J�$��n|��� ��I ���J��y��� (/�x�(w�v(/�u�(��t�/s��r�q#q�z!sK��d�*!��"��*p'+o',�+ ���f�h���n �bD�.Hs�b �J��"�*n & "GF3 & 3�����wf����3�ǁ�������J�$��n|��� ��I ���J��y����ʓ��w$b�n|��� ��I �%�J��~f����������K���H.& /���7�J�/sKdB����b���-榣�,p�1�O��cH/�F�b��#��r����� "1#>G3F3�Փ�������wb��n&�&���J������&�@�"���@?���&'�!��/���  ���F�����g$&�|���� � ��T����2H��
�
�����V�(��{(/�U���TњS2(��RT)�!���s�g"�n�bQF�b��1�"1G3FA1 3 �!�⠋��/������� 2�P���@���H��
�
� �~��##z)��3}��{�!�������� ��@��������{9����C���B"���"�)��3���@ﱱK6˛C&؉�q�|B"���Q$6��bc6���*�JQ�*Y$�Q�6�6)�˸r+cL3FG3 �f��y��3�l�<b!⨡���������9�2����2�����cb!⠰��J��� ��F������2"���"�)��3���B����2����2����̄���b

�
���(� �>(�=�HH�<�(� ��(�(�(�/�;�����v .!+�1L3G3>F3 ��&!̅�� ��	6�	Cb���(� ��(�$�H��ȩ* �ɢ�� ��ʩ*˫(� �&!̭��� �� NŽ"D�����"�I� ���bžk      �� ��  ��&�D.���b�"�ނ��J���   ? �=�. ���Kp���� 	A�� �
�)��&�>���E��� 0ދt艅E̓	E�	�W �V`�BR1����D@���TR0W�� P��uT`!L �S1R���O=E���G�TR	�S���߀G��uT	%�8N`1�W ��D@N�!��C�8T@ ޅtDN`5C��=�E�d��tTS��� 8�u�!��AT���� 8σ  D� އ���8�H�H ���D އ�� p̓A�3 ��H�H ��C ��	�T `�TS��� 0`VX�A3 �TE8LNb�GI � 0`VXCLB�$XM`	���N�/`VX� M�`�	�3R�N����S�"��T�D�H�4T@�NS���!�T@��&�.��b��.��b��.��k� ���� ��� �� ��� �� ������T@M�`	�J`G�I� �
���!�"���&����N NQ^"^�mVVb?�/��^�/�~�H}� ���J@�#d&)N7 O()~H.}�, �W�/���ne�/�#� ���D� � UL�`