����  �     	,        .   	     ?   	() 	?  T  ��������������������������������������������������������                                                                                                                                                                                                 
 @ٔ�MA    ���L �� 2��#�$3x�1 33 3XE3.;3 U  P    � �� �� �  �O����?� ��� ���5�� �                                          ���� 0  e     n             ���?���R��` ���[�[;"�o!!�{�!��=BHafI!i��I,"0�d�IJ&���a��J�IHD���!��I���a!.(��a`ia%&%F&NmbOOc���OND��N( Ai�C�D?bEi���C*"C�o�E��F��%�FNfmO&O�?�O�N�JN�(A��CDf?E&���C�*C&���E�JF�Jb(��r�� ,�!�l!I�������� ��L�pl��@>ϥ�t@	�Ft @�%%=aRc �Dt�l 	���� 9A�2P N� 4n -�K ���e;SWn �� E�pJus �խHt�c�%\�� �AP�CrR�	1G                          ��  ���&!!��(0ъ&���!���2��D�����/�P� Q�����bD﯀���R )S)�����&�&9�&�@/�D���b��D�i�ϔ�̫D����D�J S   �D *D6� ���J�
>

�堮��c��@��b���� /��@� �P? ?`��؇��� � �Qi3K&L6bMLb:C"DrA#'#[28)$)"9��1����LMD�L�LKD��������!�7�����������7��D��J��� �#�@�U���T��6S"�b�2@>�"o����""�j P F��v'�+� D. b ��l�Ub!�l!t=��!�z�<"�i;)�f��H/ 3KLf6M&��c$bD�A["L�:C���1�/�T�)��c�V� !#㨪�#Z6V� Q�j"!>W�/�Y�WQ&"Z6�c����L'"LMd����^���j_�&�Q� ���!�[I�ʪ� � 9�����4(���/�פ�ף  kq�s)p&(?���A�o �4i)3�&���2�r�� 7G� ��TTb� �YYbXYb�� �WWb�� �VVb�� ��ߛ�K ��� �$&<]&]t��� GG.
(�,)G( ,)� ����Ē�����  �@b��b(,��d�-�ś ���4��c5(�@��

�
��70(���@/�-"Ŕ������@�� &!��"���H� �̃�&!̇B�"�B!..�/���B!./�/��K �A�[)�Q�����2�(��2�/��+V"���1�/��������!�I�����%�(b�%Og� ��&�	&=�&	7��J�d�m  �����b��b��c��c��ɘt��J����   ���!333 �D�������������������D��စ�DU�RA��D	�T�`R��D�TR`�TS��� 0��@	�0T`�T@SX��C `e҃A 5�ECL�N!�G@I� `eC�LB�EM�`	�H�N��`e��M`�	�R1��N�/	�҃A5RS��P5 	�H�A3RQ���M ��L@ U4S	��4��ŠT`�a�EF��C��8� 0��TS�" R `O`�T��O��TM`	�`�GI � 0�^&����T.!�	�� @^+���E�4^&�	�G  v,�L�G�#.!��� .!�	�@Q.!��� ��.AΪ���� ����� ���� ����