����@� � @ � � @                                                                ���������                                                                                                                                                                                                                                                                                                �8�  ���      2�ӀL�G                                    ! "# $% &' )( '* �D  JHVB�� @�rB                                                   �rB�S�N  �rB�T�N  �rB�T�N��rB�� ��
� ��Ū &�����s��s�����'��᠓����9�L��0��|��7�&�	&��(��c�<(����b�a.�>�!.��?�����ɐ  �ϸ	'��"��j����c����|�9������s��s��s��s��s��s�{��� �@����0�p����� k\1��"��+R4 ��GB@ ���l��6��É����DφJ���@ `с<Љ|��DҔJ�����/�����c ���a.��?���a.��?��������r��s�!��0F����v����첂��:�<뀘��S�S� �             ��� �   �T�N  �+C�$� � �@ 8�������
w� ���4(����������c(���Ʉ���Ƀl��7�����s ��(���(/���(����/�ɢ��/�ɣ�Ʉ�ɢ��/�ʢ�����(��(�/��(���˨��'��G��&��   �����(��(� ���Ʉ�+� � � � � � � � � �    �
@��\  ��r����+�" ��&��  3�=#��2�"	�b�n��Éƛ	���/��	t�	����?              ��É��&�&'D�J�;� = ? A C E G I K M O Q S U W Y [ ] _ a c e g i k m o q s � A AA ��6� ����������Ɂ�<#a>��>"!>�6���#7�"7  ?�ך�a.�/�����`$���`.�?���#!������݂l�斁�7��,�`���f��)
.����'D.#�|􉼂�Ƀ��������@ ��8/ꁬ #w"�{������j�� D c�� �����%& +)2�������(������/����ǁĠ���t������������(d���د��Á����� �l���c���� ^�J�������J�ظ .�j��,� ��J���ЁL�0����/������ �k �(/��6 >�l�6�&ؑ�RYDښFAA bo	1�6"݀6    �2*� +0�/�������/����(��(/���6��ɟ6a.�/��!�b������!b!�|��rg$�{���������9  �f�b(��H�����2n�2X���cD���>X����z��N� � a��b�j.b�@/�n.d�ګ �Q�D�UAA bc���%&  �2>+� ������ �� �� � �W��%�������J�bK�j�J&�K&�J�W�KZ WZ"�@?�W��>����������+ ��@F��4A@g@AD��� ��@F@@6@A&��4B�nC�nDEf�F&@�9c�O��O��O��O��O� @�»(��W')���W"'ӛ�t� ['d�'��E��
` =e�C�JBFD��BET@�2ȡ�@�2���@@4�A'A�KD�JEBD�E����B@T��������ɟ������Jb@Xb!��AXbY .BBd��@@4AAt�[�\ .PPb K�O\b�N&N!.�Q&� �M�/�Ͳ��/؂����W�B@�nA�bB�nBB&B ?遮A�/�A�!��B'@�J�7�
C�b�z �Y$h4 �T�O�c��D&�@&�A&B�bC�bE�hD�J�A'ABD@@4 ��B�/�B��A'ACD���D�/���E�JD�/���AA&A�2(����/A�J W����AAt�J�XY"@�bAKb[\"B[b\ .CXbY .DDd�Y�\�"D�j��2���A�"���A�"!����'������	a>�/�	�a� ������-P��0@.��C�%���@�@@cF@�D��EAbFBbGCbHMfH�J�F�FMb(��F�2H��F�~M�j�F'�A�A�k�G�G�nFF&EG#IIc�FM�"H��F�r���H��F�r���FIs

��M���@�bA�bB@c(����/�@�@AGABD�� (����C�(O�鲠����6� �����������V5���C�  ��O
P����C��[�\�/� �����K�����[�[Kd�J�@�bAXbY .B�j@@4AAtB�J[!.X.LLb@��!����/���@@b�A&[\"KO&O .KP&P .�N&PQ&@�JLH/� �D�kِ�M�/�A��٨�AdN�NQQ&� ���4RNbSObTPbUQbVMfVO٠�SS&U�KM�/٠�U�k��f�e6���OCb� 64�T�TTcMR+S�2H��S~���S�{!S�H��S�{�S'��`��^&�_&��?���]]c���ݾ�ھ�Ӿ�־�Ҿ�ܾ� ]]�I���]^bA�k`�/�`��K&Z[f\�iKZ ]@&ABfC@c� ������������������� �BCD@�JA�J�������������}��
 BHV�W�bX ��C
�e�oF]c�������1����?��6��$� �	�F�C!.[�/�[�F�/�B������)]�J���� �A�/�A���)�Z������*F�/������F�I������]�]�9��oQ�S�U�W p�ݸ0� �*Z�����)� ��\�H��\�iÀ���:������c�����g�.�,p  $0 �*p�����u [ C�Co�C���� ^^_D��� KK�B���                    	         	  ! $'      $( 26     % 05 @E    $0 6B HT   ! (5 BI Vc   $ 2@ HV dr  	 ' 6E Tc r� �� ���0�                                                                                                                                                                                                                                                                            ���c ���F.��Ţ��t��t���      �� ӡ ��   
ׄ= ��.CÃ= ��@D S� @�#� �N�T�D � SƓ1T ��E0  ,�+��� �� ���	-c���~��}�	-s������
�b+@>�/������
|9�	'�*'
|9*�Z�	'+H?1+���	�x����+�|{����(�r	|y(�Z�)'�*'�*�*)u+>)�?Ѡ�*6�? �++7�+����	'
|9)�Z�|�� �)+s��ÁH��+�)�Z�)�|�� �  k+ E�.���d�)-T )�,�h���@/�*���*�Z-�2���@)��)'�..7-�-�2���z-'.)w+P�('�&�-�y-�-��x�(u��� +->ظ����,,7�,��,'����������w*'-�2@-��(��(�)*U�-�v-+� �-H>-.s.�)>)�{                �
Ꙫ�d���� �� ������ǁ��-.w,)w�h�-���/�ڢ�����*'01w����*کJ�⨎�b��Ơ���\3�2����+�F+�D����Ԣ,+s!N�"�+�H�����)�?.�Z--S����,�#�~��� �    +�3��J.�����3��@.�&��� ��C^�
�������͙������4�� -(.�()�� ���������� .a.�-�a-� �)D>).s.�->-�{ @*)3)~0.3.~1-3-�{ �	�{ ������/3w2 ��@�␷�� ���&��&��&��(� ��b� `   ��J� �	c	r��D ���b��b��b��� -1.s0)s*�{         ��0�
�����v&���          |                     g P                                �����������������ZtW�����0 ?V������������� ���?f
�D���/���9�K� � �\�� ��@ �0��1�  � �����&����ȁ<��+�n�h,�i,~ F���@�� +b��� �"��h �����o��� T��Ъ��� �3�M�!��  �"�@n���SD R� E �,} ��&����	B=�3��!e'&3)(3 ,|  D. "�� �$&f%�k{���o�P�� A� D��`�����%�/z!� yi(��,yi� d�y����y���x�wy��,b}(�Ģ�o�%b��w��:�:�v��6�w�,u J��t�r�գ�x�t�7��C��t����&�@?xt��	&	�7w �(w���/w���%��wk ������Ȩ������� ��7��8c�:c��i    ��x� y	wk��Ư�tl�i �� �@,u J
�+.�/��&��6��,� F�	o	46	�6	"6`."�/x(�	(?�a��/���@�'&(�('bD)�(."@n')")n(""(@n)4"	n(F.���no	�)ww��Л   ,J.
}�� �6H>����{���&���5EM�PS�Tq$""6{)��� ? ?`��؇ �#�@� �������������s�wx�xr�wx��&�3&%4 ���&3 !&�3&&%4 !%�4�*���q)�q)3p oq)&p oq)&p B�{���  c&%f!�b$niw ��%�4&b3,f�m���	�,�-yi.wk��)� �                               Y!�l!tE����@Y ("�:�       �!��&p���/��������b(����d������J�Ă���� ��,�������p�ţJ4�� ��p�(���J.����������xy     �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �U:[y������� ����l��l���6��(������ ���J�kIU�)m��k�Uz)miU�"�wk���� ���ƫ�4��l��)���     � �!�⨺� �"44c(����i�  x	� �H �

��	&�
&~4&�	Á
Ǒ	Á
Ǒ	Á
�4�J �&� �       �S��*���v���l7�,kx �%�/x$�h���@/x$�$�"@��$%b&%f���%H.%&b&�$�J� ����%�/x&��5�������;877976�06�yw�wk �,�|  D. "
o
16
�6
/6��p.
�?�/�"b�1�1n(F.��� `1�<0�b��~/H./!./����,� F�P�����   �ԧT��]���&o���	&b5�b
�b4	b
	t4�J�=��������|>�<�w{ z	P��x�&D.F&�D�� >�(϶ � !6� 7 �'!�*�>Ǩ �� &.��4&4�#�l ?4�|# '4�O �J��� +r0����(��4b���(��<a4���0�/0 @�/B0�/�w��%�w?�f����? �5� ��0b��r��r�v���wk�hw �0�/��!p��i�ǁ��&�"�x�0�J� �3(f�'&"."(b��@3�(�'�J".� �:�?x�� `�x��C�����6w � `  jq��qЛ 6����K�w� %�s��z�|q	w ��7�	~b
�b�	�
�J���)�
 ��/��łU��U(/� �!./�/x���<� ����*�)�*��(/�@���/���/�/�x���(/w!�B2�i�0&p&�Áq�0�Jwh�w岨��oq)���4�!B�H���w�4�"44b�/���6J>�i�wz�P���!�B@?w�hw�oq)��Jw�    �  �   ���� � ���  ��P�P�(���U � �2��ڃ~�ڂ8�ڃ~�ڂ8�J.
��J
� 2 ۞k ���Ě��ų&��&۞(�ł��b�ۂF�~  ��7�J.
�~  ڞ8� ���J�"� `� ���&1�&��&��&�pb�k �!1�w �    (v9�)�l()'�9� 6��o6�~6��x�w �����(��G+ԃ&�%ߟ��U  hx�B Rg�/B5r���̓��~� �)� �F� �J
��� �f�� ~ 4�h|4��� h	x5����̲�⼊�~� �h~J
 �

�2**(/������6J>V6�w����� 6y ����9�y6#6�t� �66�9�9�{ =���x��6���xw�v�9�[� �9�6��Á�� ���a���h���w�����&&&$�&%�&&�wh����	!.�3&�&3!.B2�i�q93�Joq)���$�)%�)&�)�w{ 7|!.9�?��� 6������ݨ��8�X�ݸ�8�;!>8`><�?�ب���e<�`A�e�<�[ �	��)� �6o0�����)�ݛ 796s�6栾 �khPo_��`���De�TRm�T�r�{ن�&w�� ��ǈ�w3���P� ߉ k	h$"���%�/�r��%����s�"'fX#�$!.4#bX#�'.'4d�%�#%&' &"b���ke��h�%"&r"�����M��e�s��mM���  @ �"�c)�c()b��%".~�&"b��%%!f����!��&r�%r�$v�n�ww����4n����D� K k	\%"�,f�m���%(/�����������/�k�b�)$�"����b�%�/�m�b%"��i�%��&b�miMky_�*k_�m\��\�k\�m_��H.��b�����\��(/ߠ/����w��M�wr�wm�Mw{��/xm�\�)�b��w�    %(w����� $�dw�����@�� ����3�����4T�r %(w����sx����ځl�"&$H/�$o$ N������
�()f�%"%%b(&����(�H(�).)�i)�"a&�(��#n(�"a%��� ����J "�%#b&)bD���(b����n�"d�٢%�b&wk  �4 � �      ��/   	��v�                                     ��瘰����j���������M�zs���M�kh��k�e�)��|��e�)y��e�)v��h�(� ������� k	h�)$�&d��h�+ %���s�Ǻk ��s�� ��������k�h�)����������h�ke�mh�$ N�e��M��$$&� ��\ %H%�&.&!b!�� � �
�� ۹T ��
 �	kh��M�%�/�m�M�yhk)h.�mih�)ke�蓮��e���e���h���/�󩂲����� �%h/�F�($�!�(&���$&f%�k$�&$kih�)�k�em)h�)��ek)h�)ke�ﯙ�e�﬙�h��ke��$&d�e�)���� ���T ���H� p�w���6�_�t�H�p�U�����,~
LD`�n���o�k9r��䷊�l��� ��` `�xR�  P�vq �U �  @ � ��$�`������(/�@��$�@%�H�%�$�J%$&� �$%&&�b$ni� ��$�� �kb��k�_m)b�)�_��S���b��f��&C&~�*���J�������? c	��9�sɀ�+ c	��9&)&"&6$a.'$&'%b"(b%"b(�l��'��'� �����#�(�/���#)BD)�(.(!f%�/�s�# N'�+"a.%/�@�%�i!@/�@�&O�%&b&�$ N%�*%�k$(o&%f�&�a&� �� �������ߛ  ������԰GS � Nn+4����e�#!��ЪZ�� c	��9$$&�"f%�/$�h()&�"�&�b%%b��!��#D�s�� �$$&��� �')b ��!�k).)o�@�"&""n%�"��"."n!'d���)"b��@&�"�).��Ja&��� c	��9!$�$(ba(��&�!�b��jЀ&� �%("����"&�%�%�%("%��&�&�"�J�D��/:��4!� c	��9�(¨��%�/�خ$'��$1.'0/�!����'$&�n���K���� �  �(.�(�(�).)n"'d  䤡� !D!�&.&%b%� �  �%.�%�%�&.&n!$d  �¿���� c	��9�Ԃ��j &a&�%�a%�� �)a.)n(a.(�k @"!"!n)&"&n(%"%�k �@T�� ""'6�"�(�h")6� �%(/&(/!�/�ڮ% /�&�����ڪ!�k4 �c���'�$)b&(b%�d��� c	��6$�'�%���x&�'��L� ���K�������k��� "�Ʋ�!�%@n(%"��% n!!&�%��U�p$�$�i�$���� �   ����                                                                                                                                                                 R��� L��]���� P��� �  	� ������£�   c �� �� `��� ��                                                                                                                                                                                                