����   @                                                                                                                                                                             8��������  +.  2	2'<"   +.(  "25;46"(.1  32>(+10>(#:/>(+.-0>(#.:://.:  ', 
      /+0/'*	/   : S*(*6  >#>   >$;;	:2>>6>639  T �i �9"`8�      ��/���}5�~U �             �? ������������� v� �I�C
-DHcDd @   ������ �  �/R1c � �3�2��g�Z0Y\ X        NQ Q   �9�9.#:9$ :c+ B	@ � Nt N qJ�p�,!����n�Á��E����b�Rb��l=��>�     P���B& /������>�� ���QiF��+&X&�Á��JS�&Y /�������>� P���AUb��fY�,>�   K���(/O��&V&T	&)&(?0	'�J ?�0�	0r	�z1�	�	�|(?�&�c��J�� 5�m� ��* ��b��b	b����/��t�h&��2b	�h�/�'���s-b phs&( &p-� bsph`/������( &s&p���k �	(?�/� ��%�*%/�c�������z # (��;;b<H/���;�"���;�"� ���
.b
g�J
&�ɳ�@�a�#'��+�/"�/`� ���b�b��b ���	&	(?�����ݴ��&� /�c(�'��b
�޴�?"c�� /�?"�r�r�@�{ �H���Jܴ+ ��b�C�II���̂l�Aɀ~ MB��~ PNѴ �� ��D���
 0 ����]0    ��bPF�a�7� �O(/i �Ny��m�L#� ٔC ��/�t��&�&��b��h�C�� H	*�& � 	&
&?�c�����鄠%�	%r
rs!b phs&! &pꄘ�� # ��bG��!.�"b��J��""�&��6��&����h� �,�&!�&�.�o�0��� ����ӫ~ @       )V'"W	'
r6���@&(?�6���� �������>���c��洁<�禮�7�r8�r3�r5%r4%r6)r!�k46w8%r3%r5%r7(r!�k�����1��  �   � &�&�& ��6���5&��� ��̃�e@���=��b

�
���(� �e <e <�(� ��(�(�(�/�;�����u .!��&��:�&���V��b	)bc	t�����1�	�	�r���Š*�����à*����b�%�����cG����G�������(%�(L �(��&!̹��������_�3��3�!6�!..X.��h����- !!�@,���h1�Zr��  ���>�+ ���Kr���� 	A�� �
��)��&�?���E��� 0� 0FL�`        �8Մ3@ɏ�T5V�C`!R�� @�T� E����C@ɏ�T5V�C`!� 5��CU�!A �TL ���8�	1�8VC`�3� @��
�T����>       �T@D�      ���D1� �    � N��TO�#� �8D�	�3���R1��R1R���C4*��R@*�P�  ��
N ��-+Nr�N`!NB�T��C�4��TO�# �� N��TO�#� �	� SQINA �P��CTO�A3NR`,n*��*���  1��5��91�5ͷ9�1��5��91�5ͷ9�1��5��91�5ͷ9�1��5��91�5ͷ9�1��5��91�5ͷ9ފ        "�x���"��� �" x" �$�� ��<� ���<�  �"&x���������r '�1$ �0�$��  � ��������������"�x� �"��  �"�x���"��$���x� �� "���� ���� R��������"�X��� "�� �O                                                                                                                              "�y� �*�/"�p �o��$� ��� �<8� ��� D"�x� �"�x�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        0��υ   �&�&�Á�D������(���(/������� �f�"@O�����n(/��"F��� ���)��)� ��&� ����F���Ál� >��b�8p� ?��"�����'ۼJ���F��˼ 0\� \ސ \���$[� �[���[��@(-:�00�:�� �������