��� L �C �@                                                                                                                                                                                                                                                                                                                                                                                    ������G����&��0�������?嘊ߨ?�����0�d��0��d��6�B���������/���䖔�DV�	��� 5��CU� A����?���� �����c��b� �f������K��0���D� �         �N��{������ �T� I_ � �v��_�d�����@ ���d��(�����(���   

�
�� � (���� ��)��K ���6��B�����(� ��(��������꜋ ���/������(� �   &!����� ����(/�����������(��(��B������ ���D�H� ��ڋ ������ ����������� � �� ޅ���?  ������i��J��9� � ������&��?����������9��c(��v�(?��'��9� ���'� /�&� ���&��&��@V�{&��'���T� ER���I� ��!.�6@.�/���"�k ���/ `B��0`B�D��F@�o��V�?��FGG��`�����P � ��˅�W��&��˵�r��j��bF�����rJ
��൵7��D��D��&��J����������i� � ���T���    ���������D����� ���'��)
����?����0H� ��0�kῊ&��<A(�
���K��IU�V0�U ����P ��/����/��������c(���d�&b�&����J� � ���c(���d��4�ib!�����)������(���H����� ��f� �(���H/��@������"À���)� �T5Ӌ��D   �m�mm� �	�ߛ ��䴀�J����? �BIS��@p�V���P�ϟTT Q��Q 0����T� E�S(A-�3 ��ԟX��4� 5XS �[ ���r��r��r��{ ���d��6��C��d���    �
���ɐ�TX��C � ��b��o� ��EVC`���4 ��� ��`A����$��4 ���ӛVZ������U�U� U��_B�D ����� � �������Ɩ��f��f�����H��h��h��h�����b��h����!.��"��h(��!����d�Ө!����dšJѨ/�ʢ ���������� �       �	���� �      ��É��� � (��������3 �             ��<����ʵ�T���  ���I�cd ����(?�P����L�S	� 0�P>��������㨪���ɇC ��P����GE��4���P�����`A���  �/���H�����( ��P>���P�	SQ@����?΀� �	�!>P�����d	����5��K �l�<� ���c����9� � @/��+� ȾR�IGw�JGF�t�H� �	�/���(��k� ���n	&��&�	É�� ��/�������+  �����(���������(����/�������(�������(/���� ��!��&��0�'
>��.�k���c��~�0����nD.&���^	��_\���U������V�%��e}ޗD���Shl��bU ����b��f�(?�@��/�����j���(/����؞��d�ϢD�������      ��b
�グ�� � ��)� ���b�����(� � ���)�Ș��)Ⱦ� ���� �� �������0�&�A���/�� ����)� ���É�ˠ��������c@�␽�� ���b�T��@�0� �����2(����&��6��)�� ���)��)���   ��&�� U@d�D �@��D�A��  �@ �S3 QP�4@S  @            �/��������� � ����2�@2����6C5� � S���1��5���=H@=Ȁ=��=� � TF�pb P�D��P�?y ��r��r��r��|��<��/������NΓS�`S��  ���Nԓ�Se`2D  ���BD�΃T�# � ���y@�����(��������(���@�����蟰���D�R�C� @� ������H/��"�՛�2���� � y �0P�b�L ~  ߀SY.t�J�-�)
 
6
 �(����b��&��2����.��b��&��"��i�� ���/���H�6��/����� 0�������� ��&��i�i���?������)�9�/���/���虠���������9��DD�J䀛��J�BK� �"޺ ź �h���V�y� ��
�� � �`0@�c� ����/�����M`Tă`���`��"�8��8ŀD���M�`HŀD��� ��&��?��"�c�&�&�&� � ���)��)��)� �
>�໻bF���i(O�����K���K �	!@����K�?�껷2X���b�Xl?p����P���� dD����D �	��&>�������ƀ������ ���6�O�����)� � ���(��ՠn�J.
��&��"�������)��"��e�����D�k �	�/����b�� ����)��)��� � ���bg��J� ���&��bc�����J������o  ��cG�u�� �h�e�b�                                                                                                                                                                                                @V ��D " D "� )5 �
� NP�5�8L�ņ8L���8L�E�8L���������������8\q�	�3q�^   ^B؁    �NP�5�3   �N �      ^ R�r\                                 P                                                                                                                                                                                                         