����@ HB    6'���������                                                                                                                                                                                                                                                                                                                                                                       ����������������ɀ�������h��������� ��ޖ����|�򗤘� ���)^ �
�.��l��Ɉ� �
����ݳ(�����#��ǉ����D�����'��B܃|� ����  p�ѻ �^�    ��B(��W9$�� �? �� `_Df ��QD�^D��Հ�M��_ �	��r!���6��C��/�������_��!�⹲J��c��&��0��bF�����u�꣸�b��f�����b��z��g��    �� �   ���2��b��r��&�7��2��d�2��r��&��y� �����`���킜���p�׻  9E7�O)�_�4�KP��W@�OuTBU݀U ���㉨���&��&��Ɉ�6���&��(��Ɉ�� �� ���b��"��c��t֝J��&� �թK�_�����s��{ ������������7��{�O�ﳠ��� N� �˃��˻��˃�� �� �    ��' ��tׁ�� �/�i	a>R.>*D�E��D��E��9d���7�O6� ���&�.��c��7ݨ?���X���{ ���6��2�����C��/���������� �(����c��d��#�����DܬJ��&� ���6��Ɉ� ���2�����2(���/����&��0ר/�ٴ��J� � ��� `      �'�����nM%���H_4h^�7�OW�F
aA f�4�Q�F ���c��c���J����6��&��B����s��t� ���6��2�����"���!.��&�"��c�F���&��Ɉ� ���0�/����J� ���B��r��ǉ��                                     � I� �    ����̿�����/7�O� 
��Y���T��� �rsw03wHqw`s�rT����u�r��p��r��u ���*�?!�����!.���ט������)�+ / ����	�"	`O�(�� ��&	!.�b �d!.
�b��b	�k ��
�� � ���+I��4N (L���2- �      ��������������@�X�KBx �� �  ���C  �  �  �  ��,��q  ��K �� �  ���M�   �  �  �����s  ��K �� �  �� L  �  �  �  �0�l� ���K �� �  ��`L  �  �  �  �1�l�B ���K �� �  ���@  �  �  �  �0��C ���K;
��M� ]� �� �  � 5  �  �  �  �� �� ����  � ̄r X  �  �  � ��<��K �� �  ��   �  �  �  �T� �� ����  � �  H  �  �  � �P @��K �� �  ���L�   �  �  �����s  ��K �� �  ��5L ���� �M�_.	 �� �  ��sE  �  �  �  ����Ā ����  � ��p   �  �  � � l��K �� �  ��rU  �  �  �  ����Ī ����  � ��s X  �  �  � ��<��K �� �  �� N  �  �  �  ��,�ı  ��K҃T� E� r	<? ]���@ ހ ��                                                                                                                                                                                                 ���v&xş    ���G �                      �                        �t�C ���0���7�@ �0 ���� ��dǧ�X�B�� � �XM�օ�  � ��8 `���BQ *�����_�.��k�ޠ r���? � 
 D �$F�`��~)�}�|&���{��ziy);ٷ{o�����w� �xw� ���<v.��2�����k �F���� �Ŷ�u���� �t0 v��K �&� �sΘ�̪�ŋ��K �@������+ �@������+rŔ Q�X�`7TB(� 0r���OB�r9# v��P���?�k�����������X0��� 0 �/q}��v�q ��
>

�����p���L� �u(�o�uovb��(����/��~��n~)�~)ml� n~)�~)p��"�k����B3R�8G  x����� 5`���PŃ��I	�� @x���o��R1��D�8S�nx ���'��D����$+w� ���� 6@�� �}� *��*�h� �kj)i��� �h��ji���� hi���	�h��ji����	h��� s	���*�/wg��&��&s���Ĥ�r��N�TA" �0MN0 ��0�x   ��&i��� �h*������'i��� �h*����i���	�h���	&�
&��&	
7��Ji���	�h���� �� �  ���?�����d��yށ �fr�`��`6NR�NAD�E3��`Q�`VX(�4�T��C�r�`�N0RM�`P��E8�8I, r	�N�Ճ��H`2l0� ���`@� �8ƅ1�r��(�U3�� `�S� NA��Ec��;r��	�#�B�XC�`�T��T0D�`��DE,! r	�� U`�8Y	N���R	 rYS(T "`� PT5R�RA҃b�;� ��e��� $d�&*�/��"�{ �	e����d�c��d�B��&*�/Ȼ��{��: �	/�&�c)w��b@./�/a/��/&��� �h����`���+�/�s��w�/'��&��� �hʻJZ�b+�� �� S _	������g�� osI^�/�g�O�����w ��c�(O�������J�6����r��� 1��TO�#�8�  x ���(� ���&�(���/�e� � ����&]0|�/��t]0��/��\���"t�'e@�@�����b\���"�{ 8  `�������� ����  � "|& [iy��qO�}O2v�sO�O�O�eO�kO��O�mO� @b��/��~�t�n�~��~p��~)��](/�Z�.b���Y~).�/�X��~.����W~)[y���r��}2� .�/�Y�~���](/�Z�.b����.����Y~)p��V~) Gp��Zrpi~)(?U~���,��� �+�gs�T���&+b]�a�F�D�a��j�g�+ /b� �S��S����"��b����D.X���i��
     R�� ����&��&Êl�    R�&�&���&�"�l6
.u��n�$6$"%%c�%�%.�� �&&� ���&��J��J� ����� ��� ���P� �	(y)������������������    Q� ��e��@ d�&*�/��"vs���*��w�P(���D.F.+b���O ���e��?�d��b!����!.��y�r���� �`1��SE`�	E� 0x ��n+si�@.W/��+b]�a�F�&ီg��H�g�}Up� ��*� *�w�s���P�(��+b�w�N ����M)�����i�� h��&�H?����b��y��� h�r���� �N3Ճ� 0x��r����S���OB��3̀ x �mȖ"�/�Ӳ&!�π�� ��  �r���.�H�8Մ3 x i	��7h��2�����)i���7�h��>��7f9�����T�� ���ň   �s����*�/wP�(��+b���e��?�d��b!�4�y��!�����K��8L.�$N��O��R�� >m����.o����  ݈�B�-�$��Ҡ��6�����=m����ѝ�o����� ����Rc�i�󇭀 � � �� ��  �4#� wg�}Up�u �	��	h��(����	�h����+h��(����+�h*���.�l��(��ɀ� h��(���� �h�� ���0b��/�*��v��'� � ��(?�ж�*B�����7*�/��D� � � ��@� @��)�մ��&i��� �h߲��c���� �i��� �h� �Dbgl��BQ�)�@�������o *�w�`(�w-�-L �a�f��,�hK!��hK!�b!�(�����&�,&����/�-�F�,c�,�z ,,�"���,]0z�/�,�
�u�H(����$�r�`ГRTO�#� 5E eM$MN Qx{�(Jisy�F �` �S?� wr��� G"(�@�D x f	I����v`p�����{�s(�w�����g���/�ݦ��bc`���/����*�6�6�c#*f)&S�����)&#(?�#�c�##6����#���/�x���B�_�H(�((/HG�({i����r��N�Rנ3TBT%`��A��P  �   x �*�N{�)�k�����*#)B�j ��#&� �   &ƙ�q��S� &(���ii�� h%t �&(�/��''c@F☝�'(?�(����'�*r���� `[��	��D�A� 0x��r���� `[��45N�R x ��ii��� h�r���� `[N�Rנ3��TO�#�8	�$�#�4x �@VO���DE�� DJ��Ān�� 5�T@0�                        9 �?��B���;��7�       �	��ɪkɱ �      b?�kY�qM�z>��N��ʣ          � �� ��  � �  �� �ň � �� �  �� ���Ĉ� ��� ��  � �� �  �� �  �� ���Ɉ�Έ � �� �� � �� ���̈� ��� ���ψ� ��� ���و � �� �Ɉ�و � �� �  �� ��  � �� �  ���Έ � �Ĉ � �� ��  � ��  � �� ��  � �� �� �  �� �� �  �����             � �� �Ĉ� ��� ���Έ � �� �  �� ��  � �� �  �� �  �� ��  S�F�W� �	�� �� ���?�(�y������� �      Q��r���� FP����LX� x %Ȫ�r���� `[� 5�.N�R x *�w�_�b�����'� ���FD�*.��|� ���DD�*.��ˀr���� ��OB�3RQ x E�D��򛅔TF` ���� �	*F.����{ �	*F.�!�� �f*������'� ��e��@ (d��&*�/��"�{ f	s(�����s��/w��*�/�"�e��@ d�n&�"*b����"b���r�{�"c�r�{r��L#� �Q x+�� �� �   �����? �,� 2�Q�� ��^ h����
 f	e��@�d��*bD��&7�r���� 5`U��HA�M�`��Ճ4@x f	I�� ���4(��!�_��D.����g�!.���� �z��{��� �             9	�G��Ly�Ty�?��Y��^���� ���������9&����Y��i �y �f��6� 0            � 0� �e���� d��*b����'� ��e��� �d�&@>v�/d*��X��'� ��I�� ��׈C �B�l"�B�e����d�ct�b�!.s�{ *�w��P�(��+b�w�b �a�� ��(�y������������������ �   Q׻ s	��/젾{s����C?*ڪ���� � ���&�.C�A~)�.�摄J� �    ���B�c�!N!�c!�C�/�!�����B� �*�/w`�/+b�w�s�(/��� ��w�� ��%��l�l@./�/a/��/&�/�`�+b���s��w�/�{ /���~}��}i|&�}'�r���� ���@x����;T� v�ᯀC�� *�w���)�bc��)��bcw���"��{ (y�������������ϩ�ϩ �      Q�� �*�/wI�� ��*�!���{r��N�Rנ3��ă@x *�w��P��(/������� ���� ��� ���d��6��C(����&��7��D� �    ��tv� �   !�������� ���DE FL MN TU VW \] ^  �hBL�D���a����/>���bń��'��'}'�P � ���(����@�  �h����b��y@ � h� � �����   �Ȳ��K *�w�`(�w-�-L ���-�"�a�-F.-��,&�Λ��/�,��-,�zGĜ       �
�������B�(� �(/������� ������� �	��������/���&����{ �	��� ADI�MQ�VZ�_c�fk�pu�z�� � ����������   �������������ǻ�ѻ�ۻ� �   ����      ��� ���	���# �    &*.�25�9<�A �      �@R�� �� �`�pr�o�#�D@��� 0xp�r	����E��� 0xp�r �  � -�`��8Մ3����D x�pr�� 1�#�4� 5�N N΃T�# xpr��� `[�#�4L�D`��D� xpr��� `[�SA�3ǃCL V�CS! xpr�� x����R�(�M��l#���⟽D��� � >� �~����Jr � ��3��CE 8  �ǃCL V�C`!�E3�rI  ���w��w��w  � ���w��w��w��w��wp������� �� ����l�(?�����&��0�(��좠����?���H������E���֮��&�J��         P!݇B�����#Rh�6	 ����� >̀�����