����  @ @a++4'3&"'2/    _2 :  !!!
0 ?<`   : ?>( .   00=; 
" <*3'>'=<> *-';': =':!'9':!'9':!'9':!'9';'>'=>*;'8*;'>'=>.7�Prn�c��/�����/���(/��.� +��]��2(/��.� +��^~�����S�J>ҝ������Q�/�����/�>��>ٽH�}G	�	�����/�>����Hn�G
���2�����2����>�JG�>	JG�>	J��H\�G�H]�G�� �                      �M��1 �
�� N�E0��
  �;`.    � ���/     Ql#�U31�1  #��!�!��ʺ����"��"��D� @    5����  ݏ� ��� �                                     �    ���  `       e        ��2�  ��������/�%`�,D�X�X;"�o��)�)&� )I&.�<D&\Ef)&�GEB5)3)_E"Fi���\�NFEtD�J)&�NI���\!.(��\[i\-&-B&JdbKKc���KJD��J/ D=�ؚ?@f2A&��ؚ�?�1?&�@�A�JB�J-B&JdbKKc���KJD��J/ D=���?@f2A&�s�b �J��"�*n &� !.�����?�1?&�@�A�JB�K6 ���i�K)&�)I&U������ ���&)�)��0��o�&i)�&���')�D>���&i��2���L()M')����D.���&i�N2(O�'����b��b�b�b@��D����$��F&�'9��J�D���d�D� ��O0   �#��3��?�#��r������  �Mi7G&H8bIHb:?*@r=+'+X2�"),#)*$9!�� 6����HID�H�HGD��������)�&ړ�����  ����P�P�+ UUT&U�-���� �SSb����Ț R��y���R�-���� �����K ����� ��,��bYgY�J� �QF�u�7� �P(/i �Oy��m�L#���x 7GHf8I&��^,b#@�=X""H�:?$!�� �6�/�P����^�R0 !+㨪�+V6R0 M�j*!>S�/�U�SM&*V6�^����H/"HId��������j��6�M� ���)&��9�ʪ� �6 ���� b/D�!���_D"D�nD�~\WkD .D_bEF&\�NFEtD�J\!.\Wk��(?k�2��" CC.
0�5)C0 5)� �����������  �<b��b05��d�Ѣ�� ���4��c�(�@��

�
��0(���@/��"��������@�� &!��"��ʠ��?��
� �����&�!���4>>b��u������"�>!.��/�״>!.��/��K� �&��澽w �%=�X")�M��%�!�� Ԓ(��Ԡ/�%�4R""!�� �6�/���%�����)�&�������-�(]�-Kg� �������ɐ��b��b��c��c��ǀt˽J� ���   �N���ƿ��  @��6��գ�Zd��Z�d����&��K ��@� �;��o������@@���E��� 0�26 ��㎌l;�&�/��P�   �&�	&<�&	7��J�_�d  �NĀҀԀN�̀���D���D@��TR��	A�HT` R���ET`!�T@SX��C ��	�T `�TS��� 0`VX�A3 �TE8LNb�GI � 0`VXCLB�$XM`	���N�/`VX� M�`�	�3R�N����S�"��T�D�H�4T@�NS���!�T@�T�C�@C��L USA	�S�H��5�`F��E�d�8҃� ��T@S��  R`O`eՅD���T@M�`	�J`G�I� d��D���  �����T�2H�����Pb�c�k�I@i�0>=" ��}6�����������d����3i3��A��o�0i3�0����1��Dﴀ�0ꛀ�/�c�2d�1����bD����0�e2)f1)�����&�&O�&�@/�D���b��D�0i�1������������+��+����D����D�J�8   W�f   ���ݰ�������� �����������������I�+���)�����������K ����� .��d��J��d� �    �A �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ޓ�(��@����)��J   ���� ���&��'ߝ�[-)�,�o�@ �?p����p��w� q x ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    ��}oto�nm�{|� ���f��f� g��r��������i�����g��π�ܠ/����&��I������   � >��y������������M��h6�:�ew�w@�����wST� R���������6��H��h� �   ��)��9��� ��?�>��� �������)����������TN"�  �	���/���g��)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP�����w ��:fC hRT�S����wހ F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�旓�� � 5R���Jd_d�\�	\&Cv�g: hST�R���� � �� ��� �����A�����рh�����������=��E���)�H���)�K���)�N���)��������������������y������A ��LD!  ��N C�� �Q�> ���������Y�Z�k�  ������ �V[&�-�-���-[����
-)iib��� 	��O�wC�g 2 qzw��lzpQ���U��U��U��U��U�TD<D>ADD�DTSG�S%�RA��D�MN ��A�RA��� 0	����DG�S%�RA��D	�T�`R��D�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C �艅E΃�SS� T�H�4T@