����      / (0-7)?  ?       	?  ?   ?  ? ?   ?  	!    ,  	  !  	                                                                                                                                                                                                 
  �MA        @� ��Uv(5  e�Sܽ5kZD �C��C(Od��Rb�R�iUmS 3YF3/<3     8� �� ٿ    �#  F �����?� ������ �                                          ���  ��Nw[{w� p               ������ �I�&���b�b�b�bEbO�nq&Ot�v�//�,͖/,��i8�
� k�/,��OfKP&0ObtQ&,ۖ9O""=�"!����0��Q�OPD�0����/,��!iȚ���/,�
!yК��8��D�w�wk"������/,�!y�����x��y�n��{�~�dw qv=q�E/,�!y������D�z�8��z�zwb�6�4`.z�/����s���/,�!y�����/y,�!����LO&�p�/i��Ot��v/i,"�!����O0b!P�O)�O� ���O����P����O�Jt�c�%\�� �AP�CrR�	1G                     ��zwxw|�o}}�/������w�*�k⨛�8�(��eebk�/�k� e�JP&P!.Reb�64"O�c��zO oob O���?y��QPO$�^�]�e8 ���n`.]�/�]�0]�^!.]"���n]&M�fi�oiiOOb	@~Oi"�iUdׁ�|�/���x���� /��@� �P? ?`��؇5 wxwv rKh&S NS5 ��S5 &$�D(/�B����uhd���#�`h��S5  ���S�5	���S5 sO&O�0ee&}�/�O�FQZi ���|�f��������������|���|MbfMbgi ����g��ߪW6 (��ui f����D����|�o>��/�X�5	�X�5 	���!�z�<"�i;)���G ��b�Xb5 �2b�Jr�&u�/�u������t������F������?���)�//��/�,�ހc��b�&��,�,ɖ/��V�d��6��B��b�b��b@��D���O/���D�,i�-����N�/�ܚ��D�+�D���d�D� ����c�fU     �&��f��f ����2�r�� 71� ��� ��� M��n*ڞ*��*)��J�L��n*
�*�����*)YLb��n*��*)��J��*\�� ���b
�59"��59"�� ��")�")"����  ��M�&�5 9")�.���J:")� ������F�E0(��@�
�

�"ƓH(���@��Ɣ������ :"��@��� 0�H> u���j!.i�/�J�PPb ���Nji_)�Pb�Zb��b�a�7 `ico	�<d	bbdb!c⨼�j�/�j�u�/�f�g����#����J� NP�&U�J�#�   � � ���"��&����"�n��"��&��+ ���b��b��k ���b��b��k��+� �    �v �J
�
��(��H��� ����uMbh�bs�&��?�y�Fxϴ*��?����2������s����m�#�����?�Ϣ�ڣ ���"��yC&)�F0(%��$�@��A��h����#�`h���+I� �����&�!��"�� ���&��$!;�����$!<���� ���bK�/��t�&Ϡ?��K5 	L�ozww ���n�uf]')^_&ZO&ZF Peb�&9O7 P()��ji��b������U!._�/��X�/�	��@�	j2�j�lU�JU�/����ᭈ�����!�"���&����O NR_"_�mWWb?�/��_�/��H~� ���J@�#e&)O7 P()H.~�, �X�/���nf�/�#� ���D� � �[bf !	�c59a�␖��80H
�9 .��/���5���K M��f8�����O���ꘘK X5��q"��no�#���]��s�ir��r3�&��Sl�/���� .��b2�$��������//�,C�X5 9"),F��������� ��WWb� ���� �[[b���]�      [�   ����3 v������
�T􀓶LT&�p�
�b� �&!̕"���� /	,C�X5 ��b9"),)���t�&��vK�&�)�����D�/�/,�C,y1� �!^�U�n]	&v�/�L�T�np
&e8 I�&��+ XX�-�������bO�bPOcQQc��QOtP�J��������D��Bp5jcU�SM,6"%&!!.�Z� /	, �K�&��f�2"��br�&�)�/���9")���-9��D�����J� �       �u�b&֞+%��$�@��A��+��"&%��$�?�/���#�`/�/,�zi��K ���c5��0����+Z @   ��K��K �   /,��`b-,��ab-,��bb-,��cb-,��db-㛅�@	�0T`R��	A��C��0@�������M�A��������倗�S����D���စ�DU��ET`!�T@S P�KA��T��@	�0T`�T@S P	�T�@��C XLA�	 PXR�� � @��3��@��T�` M Ք3��X�D1׋M��h6-���C��ă ��$ƃ �PP 0�L? CP�  X`���� @�UDN����_R`O`eՅD��S� �C1!Q ��MA� Q� [�8S�"����C 	� HS���@P3@X                                                                                                             \g[b���H����_�� �!����y[f\9bmg&8*)g))[+)(��%B����[�J�g�g\d\�/�[�x�/�ЪH)�u�v�ӈo !���z� � b��'{j&Tr&{&jbB!���b .brd�T�(/�!�r�kn���/��r��ޜe"Zm�7~�