����   � �5 | : : : : : : : : : :  	   	   	  	       	    	  	                                                                                                                                                                                                      y�2 R                ��� � î "3?"��!!�  �                                                                  b� +$                              �70 �                  �90��ǩ2 � �����������������Ië���)�����������K ����� .��d��J��d� �    �E@ �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ޓ�(��@����)��J   ���� ���&��'� �       �@ �?p?�/=� !�  !�� ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}to�nm�{|� i_@IQe���r��������i�����g���ˀ��������d������� � � ���������y�����y��� �����Q�!@�?>="��"��"��������6��H��h� �   ��)��9��� ��?�>��� ������������������TN"�  �	���/�����)��)��Y����b��i��F��6��J� �!������2�����2�����0��{��)����單 � �` � HP���3>"  M�À��"�"=?"�  F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�f���� � 5R�� @         �� �����"� �� � �� ��� �����A������l���Ήl����������������)��"�����"�����"�����"��������������������'����� �ρl�'��6ς,� �   �E �LD  �� �C� Q�� 茀������            �   K	��� �   ��� ��
 � �� � � ���	      ����A-��	����3 ހ �$�3�̮�̀X�O=�F]̳d̖� ��ٰ�       @ ��    �G  �������8? � U�Z��@�� ��������������Ѐ�A����� ���� p                            �����}}bh�&�~�/�Z�i� �: ~bB�k�s&k") ��� '��� ���s#�����s&�+�k()" ��� 
ks&k')  ���skb) ���k() �Ԑ��+l�* ���k+) ����+k�H��s�s .(s�(#� �됁��+k�H��PP"ssb (�s()# ����l()ks&k()# ���k()ls&l()+#� ���s�k()�+�#���*��+�^n&kH.���*y�=s%@�-n����<-)yyb �4�B��+^�nkb=sk*)%@�-n����<-)yyb �O�B��+k�H��s�s .*s�*&� �g�B��+k�H��PP"ssb *�s*)& ��yBks&k*)& ���Bks&l*)k*)+&� ���Bk�skb*��+&� ���B��+k�H��K�snrrb(s�*,�!�����+k�H��PP"Ksr�r()s*),!���kF.�Ksr�r()s*),!���lF.�Ksr�r()s*)lI +,�!����+k�H��PP"Ksr�r()s*)l")l') .�l))l()k),!����+�skb*D�(l�*&� � �Bk�skb*l�W(	l))l') "�l).��+&� �/�B��+k�skb(l�*l�)l�' �"l�.��+��+�# ��G�(�+�$֞+֞+s�k()# ��b�(�+�$k�ssb*֞+l�*&� �r�B��+k�Rss-) �����+k�Sss-) �����+k�skb(^�n%iB-)n�J�-�<-)wwb �����+<�skb(^�n%iB-)n�J�+�<-) �����+k�H���s�se r_bn$ikD.6C-n��,�!�ɒ��+Q�ssber_n&$��n.6C-n��,�!���� 701��+�Ps&se r_bn$i�n�$6�C-)n�J,!�� <�+�ks&ke r�nn_bo$ikn �6�C-)�n�n昬�o�J,!��<�+�srf�n�_o&$l�n�6C"-��n.n�o�o��*�,!��8<�+�kH.���ssb.� �V���+k�H��PP"ssb.� �e���+l�ssb.� �u���+k�skb.� �����+k�q[bpqb��qq&p�Jks&[p&. ����s Np�J��9�+�ls&[n&s)n�Jk*)k))kE (k�' �"��+[�n�n<-)wwb ���n�����n��+�ns&n). ����nD.(�niғn��+�n .ssb.� ���n�D(�n���9� �H����+�s&k") ����8s&$C�-��" ����s&+"� � � ��+�slb" ����`n&$?�-n����" ����?-)��8s&k") �� ��+$�C-)�'��'��+�'�?��+B�($�C-)���O@�+�$C�-����B()���C�-���\���E@�E�O�< (�	�ԀD�+�8"s$iC-)�l�" ����(�skb" ��� J�+��+�s&" ������s�n+"� ��� ��+*�6"skb" ��� J�+�B()*��B�(���@�+�*'��'���Ȕ�+*�'ۚ+'���@�+�9�&B()*'��:��i��ޔ� �^�嶜� ���� ������+�:�&B()$C�-��9��'i�� ��+'�����+�'��$'�����+�'���+�s"i ���$���s�n+"� ���k�H+	��?s&l") �'� ��+�s"i ���$���s�n+"� ���֮F"8s&C-)k") �G� 諀�Z�	�@7��A7���@7���� �+�s&" ����$֞s&�+�" �����?�s&)l�" ��� Z�+�$֞+֞?"s(il") ��� ��+$��?�s&�+�*"� ��� ��+'����$֞+)�'͚'͚��P�+�$֞+֞F"8s&C-)k") ���+�s&l") �Е ��+B�($��+����+���+�����+$��+�C-)��8F"s.ik")l))k') *�k)l") ���+�s&" ��� Z�k��+�s&�^�ncbo$i^p&?-)p�J."� ���o��?�-n��"� ���خs&?-)" ��$ jр�E 'r����r�J�s������]���� \��w�p��fـfɔbF�t�����ѻ���k�cq&�+�qn&^o&$?�-o��.�n�J�+�s&^n&co&$^�p?b-p��.�" ����o�J��s?b-n��"� ���q����� ��+?�(��kabn$is^bo�n?-)o�J. ����n�Jan&^o&�?�-o��.� ���n������ p���V�j�������������� f�U�s
��_�k��+�cn&^o&$^�p?b-p��.�'���n��?�-o��'��� ��k�n+c�n^boBb($�^p&?-)p�J.����n�J?-)o�J���p�+�$}�F()kH.���ssb �n))�>-). ��@�x�+�$k�H��PP"ssb }bV()l)))>�-.� �X����+$�kH.���ssbZkr)��)}�F()>-). ��q�x�+�$k�H��PP"ssbZ}rV()l))�)�>-). ����x�+�$l�ssb )i}F"(>�-.� ��� �{{b ������+$�ks&sZ'�)�}V"(>�-.� ���Z�{{b ������+$�ks&sH'l &}F"(�)>�-.� �����+$�z}bV()ls&>-). ��׳x�+�k &lZ'�)�$V�}()�n�>-)n�J�l�s.i ���z�ks&. ����x�+��k�@o&@))$*�on6oH.���ssbo}rF()>-)�n�oorz.i ���o�j�/�o�����ʋ��3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3��k�cn&�+�no&$}�F())�� �ns>b-.� ���o����+��co&� �s$i)V�}()>-). ����o�JGp&� �)>�-.� ���p��n���������kcbn�n+n�o$i?}"F())�� �ns>b-.� ���o��*�ao&� �s)i>-). ����o�JGp&� �)>�-.� ���p��n���Ø���+}�(k�H��s�s)>-)�z� {&{ )�����+�C}"(k�H��s�)�s)>-)�Z�{{b �����+}�(k�H��PP"ssb)�>-)� �{ b �/����+}�(��)k�H��PP"ssb>�-��Z{6{ )�G��္�U�T  ��D�� 0�/G���T3�/G������ ����� �����+�$[�nkbo}bF())o� >b-��o Nn�J[n&ks&. ����s Nn�J��������+�}()zlbssb>�-�� {&{ )�����+�ks&s)s . )i}D"(>�-�� {&{ )�����+�ls&s)s . )i}C"D()>-)� �{{b �ҙ�� ��A�8��� @A�8�N�T  ��N�T  �+�ks&s)s . )i}F"D()>-)� �{{b � ����+l�ssbs�  �)}�FC"D()>-)� �{{b �����+l�q[bpqb��qq&p�Jls&[p&}())>�-�� {&{ )����s�spd��3����+$��)�lZ'}F"(>�-��}()>-)�z� l�s b{ b �Y����~�/��������B����+$�h�&~n&�6kH.���s)i�!.��/�s�4���LF(>�-.� ���n�����;"��j�����+�$h��~bnc�kbH��PP"s)i�!.ʨ/�s�4���LF(>�-.� ���n�����;"��j����� ��.��LPe�.�	�E�4�.�� ��.��2 ��.��8@��+�$h��~bnc�kbH��s�)�!.��/�s�Z���LF(>�-.� ���n�����;"��j� ���+�$h��~bnc�kbH��PP"s�n)Œ!����s/Z�L F()>-). ����n�O�Ţ;�&��.��ދ�C����TA��5�B N�5�0N������ ����� ����h�&~n&�6ks&�+�$��!�⨭�s  l�rLF(l�)>�-��lz&�L (>�-��z 0{{b ���s� n䈴��;"��j�����ZrF���������2�/r��������+қ��+$�?-)�ת ���6�B�����ڴ���r�r��r��r���    	��� ��   �J�&�ą����'������&B �������� �||b!s⠛��� �re !t⠰�u!.s�/�I� ������vvb� �zzb����� yy�-���� �xxb������ ���� ������� ������S �QS RU��A@�(D�T2� 0��� %	\m&C@"-m����]m&C-)m�J�<�-y�y�+ �-<�-w�w{&{�+ %	^m&B-)m�J�<�-x�x�+ �-��� �%^�mCb-m����<-)u%i^m&C-)m�J�<�-e�t�k mm.
:�3)m: 3)� ��f�g���Ƹ����ƪ��A@�0�:��o�&�)#�:�8����P� <� � ��X�'�:03)�>����Z�)� ���㓀F�J0(��@�
�

���M(���@T�)��N������� p���&!̹"���� 	B��"�.��^�&@-)��J�<�-y�,#�2U���KM��`6	I3 �UL`!��CN�!�          S	PRQ�	A� 0CN������ ����i�������A)���22��e0�&��/�2/� ���0)�D>���/i�����r1)s0)����D.���/it�1u�0����b��bYb�b@��D����$��F/�09��JZ'���௺D����D�J >u�   �/+�9B�LV�^i� �-�-���M�����GL*� 	  �@����Z'���6ȟ�k����k`.li�����K    �ib�5Ǭ6'7'�� ���n�^b�$i�� �6�?-)���D�怴J�� �ڐ��b��b��c��cٞ��t��J������]Y�^I�@4�Re��-�̀F� DT  �� �� @�  � PP��@̓0� 4 F����G�'�8"�b
�� F�������ho�����&� �F �������6��î�b��������� �� �   0# A�L	�3 � ��  ��  � Ҡ �� �� �� �� �� �� �� �� Ȯ �� �� �� �� �� č �  � �� S U @Pmh�@��NĀҀԀN�̀�D��C��T@SXGS�TR���@MN0 ���R��C 	�H��HGS�TR��AX�K@��� 0�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C C G�S%�RA��D�NS��S!�D�H�4T@                                                                                                                                                                                                