��� L B012345670123456701234567012345670123456701234567  #2. <1#21+5'=----  #2*	    ;$:$/2  _:
?5 8` ':���������                                                                                                                                                                                                                                                                �����?���� �&��J���������0��� ���k� �D��		c�	c�b�����J���bD����&�D.��!����!.��7��̠��� �        @         @      @    'ӛ�t� \'�G�O@���_��P ���&�0 ��Z
��c(O������d�����c����� �	��D�ڢ���@���/�o�zN

��&���   �
��"��b۳bܠb��j�ҪΠ���c�J
��

���J��0��d��0��K���ڶJ         	b�n���J� � ��	&�`�� �	c��	U���P@���!�ڠ/������ڶ���&���(����/����(����(��@���&����i���(���h���j����	�� �"�b� �F.��+�(/���H��b��������� /���ڨ/��� ����� ��c�(�������F������8����������� �  ��� ��0 �������� &!�ʀ�� �����X.��c(��

�
�薀8��J����o��R1��D���� N$ �[��D� �@C����	8�T5 ��&�R���D�8TT Q��P ����/a� � �f �l�瑠��z�b���D㉬��6�.D�E��p�  ?@ ��&��&���(����s�(���  ����� �������������������
�T � ��'� �ŉl�(/ŖB��bF�����&�P.��/���� �  ���� ������/��)����ȟ��"����(/�𢯁���� ����ʀ�`�P� � ��?@ ��`����_��`P�� ���b��b��k � ��l�&��������F�����rJ
��ಲ7��&��D�����������d��'��    �
   ��¿�l��0��&�?� ��i	�<bF�4.���� ����?� /���� ��¨�܃��������`��������}���� `��/�h �� �Ϡ���&��&� F���b
�������	���)����J�O���������߭J��������0��r�i��&�"ޒ�J��ޒ��������)�����&��)��)��)��J���ޠ�ޒ�/�ޔ���    ���!���o���� �8 ����v��� �oJ�g��T ��� ��&��/�����T�A 4� �E#0 �������� �  �00�00�qq�qq̲�̲��������44�44�uu�uuݶ�ݶ�������� �	  � 1��5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ ����&�����mm� �� � ����  �� ����8