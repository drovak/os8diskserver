���� � � ��> -19??->"=88?0>���������                                                                                                                                                                                                                                                                                                                                                   � ��,&BfCb!�⨎��F��'⠛��&(?�-��-'�����0��,�����/���,Xn��ޖ��&����b��k X��Ш��ϴи� �Б��V���'�.��s�{��� � ���b��d�-6��B.o./6�-�.�//--t.�J���� 0    �Ѣ��X$���x��� ���#O���!E�,!.F,d�&�-&��.cH��/.b��ϰ-������6�?-(/����l-6�6C.�l�/&��� .D.�	&/�"H5�4�h,	'�	�/!.	�{ 1fD�1F.1�1.� ��������)D�J� �5q.,,&4�!+�++b���BCf��� �!��&���^��00�0H � �pqU�X$,!.G b�!. !b�!.!"b�!."#b�!.#�i bD �,,&,.,bgw �J��ï�c��-(/����l-6�6061626.6.D..,"	�l0	'1	'2	'�"�DD�,,&,&!D.!,",,b#bDD�,,&,&�����c��-(/����h-6.636� ����!�z��"tuU�r�sXT!3�"H�//cD/�	&3.x/�/@.,,&��,�"���,.�	��	�3!.	,r	3b!�����	�/�J.�'�,�b)b(��@,�,o�,���/�,�,b�b�l(?�-��6��&-&�-�-c�ǉ-��ƪCBf���B�C�i�[%2"_l"��!���  �A�o �4i)3�&^�Cu�Qdr"qX$��"�/���b	�l-6(?�..c(��/�/5&4�lZ-ਟ�.�)�/�.5&��)�,�	�y	.r	/r	t"�J#�/���b	�l(?�./c(��./b54f�.��H.���,	'�	�.!.	/r	t#D��� <����  ���B��b<�c��K   ��'��{A�� � � ���ۀCX�A�
Z%A.5n$4&�,�+b%bq6�$�!7�&�'&�'�=&�<��-��-"���-��J��&-� -�i.�i.��8..C@�9��8F.�-�)6O79B-��6��7��� ��J>

��ʃ�ʄ��8�Bb�C������ʛ � �H/��"��� �@ �?������ �@EO�  Xc�^���A�%�q6�$�!7�-&&�'�<�F.��b�-d�����&��-�|6�J7�J��&F-"���E�"���-�J��"�o-�z��&-G".-bb	�l	?.t��� ���6.����d.�DDcBDdDC6���S�[ +F��+��� ��&�	&�-&	7-�J�?��>��"@�@����K�� X��^�4��?˦���b��b��c��G��D�(���i  p �
��&��&��4��t��J��'��'�����*� @?>f�A&���5�??&4�>H.>?b?�@.@Ad�?�4@b5�kC�iO�)�����r�*r(��بi@ @ �� �=�J��h��B��b=�b��ǁ��� � �	� � �
쭿��� �����4����q���2��|��<�������<--b
���-����-r������|��<�(V-�`-�-�-`.'�/�-�''b!����7�����s�Θ��'H.�����'����������2�����'��� ���&�	&	7��J'+&倿 �  �HP�.�/��P��5C����x���$���U�l >٣_ `����  !�������b		c�t�עe�-�ba-/������..!.H-�-.b�r�����-� �u���٢����r����'� >��y�  ��ؒ��r��r��r�b	c	�t���������������>@������&��É�ǁ����J��� i ����������  �� 8[�� �-�b.-cJ
�
��-�9-.D����������� �`  >��/@)[-"DM͚�R�RiRiRib����J
��l�0 ��#�z!�����S)S)T�����&;ӔR���R�Rik�������/�V��O�r�_�ǚW��\.x��Ot� �	X��  ��x�ꅊ�����                                                                                                                                                                                                ���&�	&��w�����	(?��������   ������|������H �
�.�ǁ���	���Á���8�<@�D �� ����F �����������F ��H
 �́��.����&��� ����'8� ���/�ڢ��tӁ�����b� 0�������߉������2�� (��i  p ��ᴐ��  p  �����0��,�����/�⢨��գ&��À�l��6��'�����t���V���~��'��7��I��/�߃��t��D�����r��w� ���� �Შ����'��'� �             �������޶j�O� ��D �������� ���qL����m�?x�����