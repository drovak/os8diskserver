����@ HD �  	  	 	       	  ?���������                                                                                                                                                                                                                                                                            ��� �������8���1�����/����.���N����?���^���Or����;��_9��n�7�~/�����,��o���w�������+�����������1���;����=��|���h�?���=����w���=����    �    - � =   M � ]   m � }   � � �   � � �   � � �   � � � 7 ���D�⢠���A.�����Ɉ  �
��B�b��b�j�����ÿ���&��0J
��
.
��������C�(���(���(/���(��@�����(/��B��L������� � �      �<�|��D��J��� �.��"� B� "� ��  @��  @��  ���  @��  H.��  @/��  H���  @���  @>��   ?� � N� � O� �  � ^� � _� �  L n�� � o� � ~�� � � � �� � ��� � �� � �� �  H���   �� �  @���  @���  H|��  �h��  ȿ��  ����  ����  ����  H �q.8/�H�&/&{�bb!���&&��a.�/��������a.�/��������&������j&&��/`i��bba���'��r���'�����n&����������66��J� �   ��ݟhԿK��G�XE�HI�.�/�>�Z.ࠖ��@)�@)��*J��@��@�����@X�>Z�.��J���"/@)���Kԟ�E��P�.�/���@X�>��@���@)G �<��EH�P.����; ��@)�<��E�HP�.�/�;�Q�"@K��G��(��𢯁���� ����� �F��  @G�� ��?@ �Ho(K�8�o��� �������&���� p	��˴������ ���2��l��� 	 Ӵ���΁�� �����  ������r��s����'��� ���h��h��h��h�o��4����D���� �   ��4ˁ���@�R�������!�ۃ�� �!��&���p��������������}��
 ��  �� �����R������� ��������D����������C�O� �����������Ĺ������������������������������ ������������?�������������������������������R�_����[������������]��������c�����g������������f����������������������� �/����?�>������ �
� �  �00�00�qq�qq̲�̲��������44�44�uu�uuݶ�ݶ�������� �	  � 1��5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ1ܳ5ͷ ����&�����mm� �� � ���� V�� ����8 �	���H� ��(� �����(��(��� ��Nr`     ��ˈ���(���(/�@��/��"����(/���˭� ��HN��6�?�
�

��(��������� �   !��&��� �     ���ڙ���x�ph `X PH @8 0(     �	���]�A   ��
? ��� ���6��<��s�F���2��s����r��g��â����8�(?��'� � ���n��b���b�� ����?����c ���F.��Ţ��t��t���      �� ӡ ��   
ׄ= ��.CÃ= ��@D S� @�#� �N�T�D � SƓ1T ��E0  ,�+��� ��X`��$�R�	C�8�8��1MT�TMN R���CXT�T%����@ ���ES� 0R��NBS�`�UE�3 �  ���UET3 �  �L`!�Mu���BC�8�P`���T�5�E3��@�v��DO�#N(��E3 I�NB���D� 0                                                                                                                                                                                                            Փ@�P �W��C �  �N�PO�#�FqRN�  � ��c`s�8RM TR�IC a�t�E��CЃRN �DU3P#��� �UE�3��BR1 �C���u�C�U�A3�8Փ@�P PR��NBO�TDQԄ��C TTTpMN �WNe �g��C GT�����Z                                                                                                                                                                                                 �5TX�R���DI�4N�!�Nr`�M�P�NBρ`W�8������C	���Cq� 1�Zr`��d�OB�I3�NB���8TTpMN �T�MAR���D� Љd�8ɇCY��X0 ���CX�SA��C	���FaN`!�EES� 0I�4T� D�D�2��Dd��������D��� ���޴                                                                                                                                                                                                ԉD�	8��7C� �M�P��G�d�OB��4�X0���	8�S5R�ND!���	5� 0۠3�EES�8ٔCXR��AT` S2 �W��T�5                                                                           ��:^���������                                                                                                                                                                                                ���v  ( �����O � �                   ������                           O � �8ɺ� �8�׃����  q��͌�L� �TY<�4E�� � -���w� a               ֩AR?�(�i�s�
��� �v���؇?����� ���  �&���&��ff�$&�%�#c�(/�~��b�(/�}�@�␪��"P|���#{"���#H.$ &z ����                                                                         z (��~z ~)���R?�y	� 
���wv{B��; �2bb�b6b�b�b�l���t���;	���ɼ���� ���b%b��?��2>IZ\�+]b,8h$2t%'�¨�����Ai����Bɚ�/�D�Ր�ʉ��< ���� ��Á��@���<�����@)G<�>����"@G�u@ee�@ BPl����K�O� ��$�����L��.������&M������X�Ni����K��������&N���0(��@���Xn!.7�Bt'�K��G�� ��/���@.��/�;�HL�N����>���/�R�Ri�Ri�@)�7�@��F�@)d�@�X$�t%'��6Zi!.7�/G;�H  \ t��8��z  ��XI�F��\Xi�\��X��Ԩ�&f�Kܟ�X�.Kiإ�L��D.�����$�;�%H$�����"H��Q)M�����"!2���ہL\�ipO���28(�|R8�2t�.��|KԟG�� !���ہL�`��{��+��D. b ��p�Yb!�l!tE��!�zD�i�)�@�ZL���1f.���>��&L��hࠫ�N�Q�Q�Q1�M�����\1b!���i O	���;�H;
&1"�&8X�r2d�9��9b�9r�F�@)2@)0&1 .1b!1�1�*�R�b�R��R��l'"
��JX�
X~$
'%
'��0bKië�EH�P��k �88�0�uO6�<�|1D���@�X$�22t%2'��bZiGV�����K��G��W�G ��\b!\� �� ��6�)B!q�0/�;�7�;)�b�&� ��96�����9B�8x'�&��8��Jr�9b�g���<�XE�HI�.>).�/��"@Z�.��J���"/@)KԟGܺ�*� �XQ��[��xO(�<L������N�7Ki����&�&D�B���A�=V�����=i��J�ܖ�@)�2&B��ݲ�b�i�x���6X�$'%'X����@)�� F2�@�@ے@7��@)7Q)�Q)�Q)Q)BZi6&H����b� �    ����� � ��@L������;0�Z�N�@H�`� 8���F���f<E�HB��F��Bi���bc(���c�/�E�H��&�?���FA�=ߓ�?����@)@)GD�=T���;=�H��F>��U�(?�ʦ2��������&<��ˡ�   2Ki���EH�2�/�B���� ����P.��;�G�3�b@˛3�/���@3����0B��!@������A��
������[] ��d��4��b98h��6��C��b(����	&��&�	�a���?�䤘��ƛ9&��K����&�9&�d���"��h ��Ǜ'8���~��&���r9�b	�l	�<�tǁ�� �a.���ϘO϶���&��&�d�;�P       ����(���/���歿���� �����x[� \F\�D\�]\&F.�� `��)3U).U)NU)�R��b\&��@����,��<b�|��[�������&�\"�����b�l(?�!�\$���D�J�!�l�\�t��*��&��*<���Ki���KI�����D�E�HP�.�/�;�\�@�G,�<L�\ ��|�EK�ksW# �"`�!@�I� 0 Q)&�Q)Q�Ȥ�B��(/��� ���Q)������E��Kן��;f��U�L��N�Ti��� ��S�S��B���� ��B����/�(/U���bc(��c�/�R�(��c!����Q)Q)��F͚U�FR� ��R�Rik;m�� � ��(0 l
�*4 � �^Rf�������T���Q�Q�Q�R�QE��I�Z.ਢ�JT��.�>��/@)[-"DM͚�R�RiRiRib����J
��l�0 ��#�z!�����S)S)T�����&; �R���R�Rik�������/�V��O����ǚW�� ��O� �	X��0 l'y����� �f� ��/���;�	� �Ti���\Oi�����/�P�8���X.��/�Z���.�>h��@��8�.6��.�/�>�\@/È�@[�.'X~.-�Z�9� F��@��� E	�P�.�/�;�H ����@)�+ �3�k<�����@K��G�� ��@)R7��P�H���4K� �8 R�e `?����&�6�6>)d�bc�c��b��[ ���Z�ਥ�J����I.[ ����>)��2@��Z�.��J��.B���� �/�/@)X.���/��.�/�[�'�{��/��� w��2�;�#�6T��P�.�/�خb��b����b��V��&�ך� �   �>o������ B	���P��0��8U�� �B���@.�/�OU�� Y��(��]]bD�⸖d�&\Yi�^��_&]D.]\b\�_�J]^"]d�O� ��X� ���&8�'�9��F�k8�rg�;�4� ����֋ �!��&����<E�HP�.�/;\��@)G ���Ѐ��?�8 ���
�� �&���k ����k�C� ��&�&� ��&�&� ��J����(/�� ��(���@.�/��"��K ��n&��; �"ȼ�;G� ��r�/�º B	���(�� ��(���U�� �I.�>.�[��Z�.��J���"/@)� �             �I�����a��� ���\FO������\FO	����� � �"b8�� ē�� !�&8(�|!�K� ��2��F�[0���X����s���>��@)�$��{  � �d������Ë����Ë; �� �dn&	&	H?�[�����/��"	@9���@)� �  �`(� �� �            ��A \]f^_fe�fB��� �Yi�d�]�"Ș��/e�J�Iabfdc&����/�B��������JU����B����/���B��� �������!.U��b\�i�/!.e"@��!���*�b	�b��	c`	ca	cb	ccb(��H/���ߚ򋒠����K�彠��π�����# 
�����<$� \`�&]�&^�&_�&��&]^f_�i�H.��b��.�o�鄏��\�h� �      ](/^(/_�/�ڮ] /�^�(_�������\�\�j\�k ��fn�@n��q����Υdľ�   _�/�^��]�]�/�_�� �@c�__&b�^^&a�]]&� ��       �1��-��f�fff _
ܯ Y��cbDD�D.c�* ]H]�^.^_b_�\�K� �_D._^b^�].]�k �(�� ��U�� �Kޟ���\�b�b�hG�&���x��bF�����rJ
���7�JB՚��/�;�ZH�"� � C	կ� ��Cؚ��/�U����\�K �}������  @�N�"P� �)\P� X��\Yi��]Bi��� ��X�Bi�����/Z(�U��d�A�\F.�]Xi�]�]Xi�^�]�"����&��(��]�/��^�/�����&���J�DɈ^�� ������2Ӂl���  ���ɔɹ�������  � ���   ]a^bb_bc�i������X�Y ���� ��r����BH�U<�XE�HK�Õ�EH���c�d��F)G;�gH<��XE�HI�.�/�>�Z.࠹��@)�/"@K��G��X�>Z�.��J���"�J��@)��*<>�EH�P.�����@)A=����D�=T�����&?��"@�@K����@�G;�(H;   ҏ� � X� 0��� �U :!�� @+ 	_K�M������ � ��@փ@� 4֌@� 1֒@ Pց@��@ց0��@F�P��@�P� 4��   �&�&&�J
�
���9D�������!������3G  Ϗ�TC � ��4E 0�� ���LR � X� 0Œ E�!Ɓ� @�� � ��0� 0�� ��DÏ�T0 � D� @����������� ��Á������&��Á�π��D������c����l։<�t���	�(����n���   ��.�ǁ�ʁ����� ������w�|������ ��Ȳ��r&�b��{����
����� L��]���� P��� �  	� ������£� .���J8�����������  � ��%d$� �䐖���&��&��,��|��K ;������  �����K; � � �૨� �T����Zn����D!���b�&
&PX�.[w
7��J��;   B՚�(?͠OU͔��� ���?�>���<�?�>��@)@)G;�
H+� � ��� �� �  
�� � ���F�@?��OB����4���� ��@)��?���,�c+;c����@�  ���"���;1���'��'��Á(����� �   �� -���-�/��"@X�--&� �Kԟ�E��P�.�/�;��"@ś������   ��� D���C���à 
�
�
  ���Xq���������χQ�����l� ���F��4��bd(?���(��������#��n>��@�@؞&�� � " .�   d&	&	.6	/6.� �kX����_�֏��_r�o�گ  � �� �@ �2�/�\��@)]@)� � 3�             DT  �� � PP��@̓0� 48C �@`}��]�&��(��&c���&�'�Ö�j��Á�����ʺ������7��DҜJ��<��Z
��ǖ�'��7�(6�*6�<�&|�
&�	&�X�
	t��	
g	�J�����r��{&;�=!,��  @ ��ٍ �� �� �� Ҡ �� �� �� �� �� �� Ԁ�������߄������ ����������0(��H
��桁��.�ࡐ&��� ���'8� ���/�����t������'�l��0 ���>���'�"(����,! �'h/�!�''&��'�'�!�����������\Zn]Oi�������b
�l�<�(O�
�f����6�.�l�<�
G�JO� �
��� � 0�[ �����O ����8�<���Ai=b���EݚP.�����@)Kԟ��DE�2Bi���(����/�ᢠ���@)E�~�E��G�UA�=Z�����EiHP�.�/�;�	HKן���D�=n�����D�EH�Pᒨ��.�/���@X�.F�@)�2��G��@)G;�DH+   ������� �� �       ����� �E� 
��P�@��pK�                                                                                                                                                                                                