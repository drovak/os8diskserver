����  ��� 	   	  	  	    	    	  	 	  	 	   8 	     7                                                                                                                                                                                                 
 9"`8�    @�   k^�Ѝ̀����'�������i � ������
��۪�Ǫ�� �� I�6�+� @�P �      �  F  � ���?�U�Z �� ���� �������                                  �	'   ��
�Ĭ��o � !�������}��o�oP"�Qb�:�U;'<'��<9��9�D8�Z�ndb8()$"����d+i$�� ���
8"('��+�'� ��8"(��!˚+��!����8()�!� �� ZFBo8"(?��*i�x�&��d$i"���+�d$i"� ϐ	��
 �� �i�6)��
 �� � ��A�]���i�6)����  ��i������� ��]�^]bi^b.��^��]�]�/�^�z�/�� ��6�N]&�^�^i&])I��]�]�n]�/�^����^�j �/�]^f]i&^)e�e����^"^o]]B���^z"��� �J�瀱��cH/�F�b��#��r���"���2Jam�ԃR]&^�_�`�a�I�Hp&_i&^)��ai&`)��p�J]�J �� Z�o��9�����9����+�qd&�9�]�n9^&^D.()$"����+^�]�J ����+��9�]�n9^&;q"d^bD�C()*$�"���+�qd&$"�����+�d$i���^]D�� ȑ�� F.b�7� �P(/i �O �Z6B
]&�+��;�d�nC8"(]�*��$�"�����+i�()���d�$"����8()d$i"���]��� ���� �	Li&A���iiA�* �4�*L"iiQ�*"iiQ�* �B�*R]&J)Li&]O 38r43sr���i&]O r��J����]��� R�����6)�˸rc(��6��R]&K)Di&]O 38r43s����i]bO	��*K)���]�J ���*J)84'3Lri&���+��ii��*J) ���*K)84'3Lrii��*+�"ii��*K) ���*J)84'3Lri&��+��i&��J�� В�� �8�(�/�;�����v .!��&��:�&�4�R]&J)]O 38r4Lri3c$��]��R�]ii&]O $��J����]���  ��R�]Kb]�O384'Di&39H�:]�JR]&i�]O H��K����]��� %��R�]Jb��84'�L�i]bO533sn�����i]bO5n��J����]��� I��𫀀1 �
�)��&�>���E��� 0R]&K)�8�4�~Di&]O 53'39��:��i]bO5���K����]��� ���R�]Kb]�O53�~84'�L�i3cΓ�]��R�]i��i]bO5Γ�K����]��� ���R�]Jb��]O 53'�8�4�~Di&39��:]�JR]&��i]bO5���J����]��� ϓ�o�8_&R�]LbiOb$��+�x�&]H.�D�_"(7�)]�O*	E^&$D����^�J'���]��� ����R]&iObJ��+�x�&]H.�D�_()7))]O *E�^df$���^��'��]��� %��G�]�n+�Li&]N m���i]bN	m�Jy�&�+�cdf,#����]�J �K�L�� @         U��@� G]&�+�J)Li&]N G)��Ji&]N G)��Jy�&�+�rc&sd&,#����]�J ���LR]&K)�8�4]rO53�~Li&39��J]�JR]&J)]O 38r4Lri3c��]��R�]i��i]bO5��K����]��R�]ii&]O ��J����]��� �����  P����$���
�`S�R]&K)�]�O384'Di&39I�Z]�JR]&J)�8�4]rO53�~Di&39I�Z]�JR]&i�]O I��K����]��R�]i�i�]O 5)I�ZJ)���]�J � �Z�+�f����o8"D()�D�d6b*؞-�-�-'��$�"� J��諀�Z�|�A3"p>b'h���X Z���  �@���+�7�)o�8L"(*��-�-�;�-'����+؞	d&7))o8"()*'��$�"� �����+J�3�84'8o"Li&7k&�d�3j67�-i�-3�=���g�gD"������3�Zi4E4H>���3z2��� ���Z� �>')h)���%�|p&i)�Е ��%=�"��%����%���%�����]bo8"i�b?�|7bk�n{i]j&7�-i�-]�-���g�gD"����d�g	 ���x�&�{�����wҿJb���]��i�i: ���]z"��� � �j�{�]^f8"oi&7))i()]*)'Κ$D����]�Ji^D^�/�]�z�/��J)�w�x��o �@�j퀶 J���긬������	�w��H�����{�]^f8o"i7b)i�(]�*'��$�D�/�]��i�^^B���]z"����J���w/x�&�� ���F�ai_n``bi_b���J����a��� �� HaiNGpi]n^i_n`Jb`�84'_3'^i&])��j`D"i_b���^�i]b���`�i_b���J����p��a��� ����� ��Ha&]�^�J)^8"4]r3y)�z^D"i]b)���)�z^i&]))�zJ)���a�J � �z�a&�OR`i_n^^bi_bL��`��^�i_bL��J����a��� *� �{]f^8boi&7))i()]*)'ښ$D����]�Ji^D^�/�]�z�/���J)�w�x���o �M�z���"i�#��#9�
]&�a&�`�]_&J�*`H.�R�
]"_KbG�^bfbN 3_rDG�337��84'4D2i3c��b�<b&^�J`�J�e��`�]_&�`�H��R
"]_&G^&b_bDG�f�oi�bN f)��ze�/JJ"���b�>b&^�Je`d�]�	]&a�J �� p� �nz�"�k9b'k����ip&(����whbp(i�ߗ�]���^^b@C(^�G*	'��+$����]@ C()]G *'��+�$��������9(/�D�!8⨰��8�8�j����8�2/���=���+Z�[�k��D?�8Hb[ZfJ)84'3Lriiq��84'Li&q� ��
d&x�&g")����+��iiq�J) �S ������  �J�H`DD�O�G Da9b `�__bD8�_)+�_`D�_�9 .`_b�����__B`�/����`�a�J_9b `�_)����_�`�J ����� �Ea&9 .`_f_D.8_b�^6^H>���6Q.�_���@^�^9+_�`�J_9b `�_)���_�`_"�����`ad�_�9 .`_b뚈��_`D�� ������9�'�� x& ]) �a9b `�__bD8�_)+�_`D�_�9 .`_b���x���j__B`�/����_"��c^�b=�&_D.8Kbܓ84'^3'4D2i3cZ����i6^)ZؚK)���_)a��_�9 .`_bϚ���_`D�� ���� � D(i�()�d�$'��خd$iD�/��D�E�����8����v&��	�l�����]�nZ�l]]&]? 8o�^���_o_)�]�FE���`]bFL���]i&^)�Ú�]�@4]i&^3'`�/^�ř�`����i ���_)�ê_) �����ǯ�D�?8�[�ZJb8�43wLi&���B�8()*$����8�4Lrii� ��
�dxb�gb"�����+�ii���J) �� ��� ��}6�����������퀳�d����2i2��@��o�/i2�/�����0��Dﴀ�/����/�c�1d�0����bD����/��e1)f0)�����&�&M�&�@/�D���b��D�/i�0�Ȅ���������+��+��D����D�J�8   W��f   ���ݰ���������}� (R�&����ć�������'�� �nnb!d⠑�� ��c�N!e�/�f�!d⠙�� ��R⑙f��J��J� ��R⑙f'�������������K ��ggb� �llbklb��� �jjb��� �iib��� �����K ��� ��� �X\&�-�-���-\����
-)jjb�J��$�� �-
�-h�hm&m�+ �X\&�-�-���-\����
-)iib� ��7�Sbtgt�J� �u�n7&Tt&u'u .tt�A��{քo
�������+i��(	�+� �i"(� i��i�+���   �	����$I.��)ڞ-,�&%�2��+T�� ��n8()iC"o()�*)'��뀷Ԁ�!Iu�� ��{�|6�iB�o8()7))�*)���d�$D����w�$|�{v�*g	 ����i�FE���{�jx�* A d7l&i@ !l㨻�i@ �l�l!>j�/�j��֮St&llC!d���d .dtd�l�A!.l�?�A��خd{b����{�x|'�d�lm6��K}V',)�Є�����%�������������ߗ �X\&�-�-�-�\�J�
�-f�X\&�-�-�\�J�
�-N�e�k \\.
@�)\@ �)� ���������� ��  ��Y�&�@ �)�.�枼J�)� ����ɶF�H0(��@�
�

���I(��@��)��N����@�� p&!��"����   +�r���� ������(% �r� ���6��B�8bo()�+� �΍c͍di: o8"C()�*)˚�d�R�&$D����Ed&gB"���i"(ڞd$i'��E������JЯJ�خd$iD�/�i��(	d$i���x�'�v�� �  �A���F.��b
����b��z�.��&��"��b��r=�&���H>��+ ���$                   ����}�o������Z����[}K�+退D�8� d7l&i@ !l㨧�i@ �l�l!>j�/�j��l��T�tlc!d���ldB d�t�JTt&dlc���ltD�l�!A���A�*�d�{�/��{xb|�~dlcm�d���V���&��&� 6 W0� '�D��� ��r����̪�ت徥ǽU��U�V*ffd����������������D�����TSG�S%�RA��D�MN ��A�RA��� 0	����DG�S%�RA��D	�T�`R��D�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C �艅E΃�SS� T�H�4T@E�N�Ƀ�ʆ��O��8J
��
.
���8@������/������O���&��0��&��HO��� �怀4ɀc�����&,�������������L� ����� � �ʀ&����x��h�����r

�����$ ���T���/����d����j��&�� 	�
���b�ؾ���   ��� ���R��C 	�H��HGS�TR��AX�K@��� 0�� ��A�RA��� 0G�S%�RA��D	�ɂ RA��D	�	��R�H��C C G�S%�RA��D�NS��S!�D�H�4T@� �                                                 � L B �/�¢h#�t��R1�� jfi)  �����)����F��阾J
�
��.�T-  �B���?<�����b�����(����/����(����(��@����&���ݢ�!|�ԫ�����d��6� � L �ۢ�݂��d͊���  ��������!333 @J
�
��H���                                                                                                                                                                                                