����  �$1$2=*!*  : /#/#8
8
8
"=#"=#*4  <(./<(+
=%9.=%8.= ??     !/##<(///"
//#+88  ';/#988/';/#/#/#  ##8
8
8
%<#%<%://};:	 ;5;0B A3,'>                                                                                                                                                                                                 ��i� �;`.�� � ���/�  �  �$i� @   ��    �     cj3o\3t 8 ���P��"�1#a�" 3O�!*�1X�S$3F"����LA  � �       � ���@ ���%�s?�����      ��w���8�� � ek"��"�  ��������/�%`�,D�F́3ɀ39VD3�04IT�/���3X�V3I{4I6�FU W(/�a����V6)�H�(���3��4I6F�Ua(��b�/�V�6��3����C4/��H8i�'� ��3G��49/�����3�t�BXbZ�n[4iZ�J�V�6/��c����FT"���F6)FU FFbY�/�F���Hs�b �J��" @��8#�!.�/�\�F'\�jWZ&�[����F.\[f�\�F'\[d�/��!.�/�\��zC:i;<��`2@���`r�]v��7��z���!F�TF�_���s^D!]���z=���/�7���?���`�'�5�� ����� /	3Ǔ�49/؛���/�-��b�p�   �
�@.b/�F��� K"L="J>"D� �C�ȁ�EI&�J�������IJ"�* IF�J� ���DH/��O��� �	l��En!Eb1%�E�+�J!�/�3��[�!� /&�� �f*&f�-*�c1%�.��� N������ ���*bfn-i*&19%��� N�]��ի����� �P(/i �Oy��m�L#� � B�⠇�3є�3��4I6F�Ua(��b�/�V�6��(/�3��4I6/�FU a(/��� ?�@b�Ab��l����D"ˤ ��B⽾f��̯�)A #� �       ����    $� �����FFb!�>�F!.�/+F�� ��Q�Am2��J�B�GGb��KB6)b6���A&(?�� ��  GD�Cm���J���� �,��3���34/�,%���nH1i��� 0	�(��� /�0��� /�0��� ����K ��<)D ���<)D ���<( N�Á(�J
�
.
� � ���D�/��C�kC�/�ۻ ���������=�(�(�P� !��&��<�� b �d��� �� 6� C

�
��  4��� EEU (��S /���RP" ��K6)MH/ON"6�� &!��"�Ϊ ��K�6L�6�� F6F�de���Ff h�cXh��~h.h��G&G(?��g0h'G�JV6)4��3�� 3��499��3���49�9�3ɨ�3灬3����:3_��@���E��� 0iV�q�� 5�C�`CAN2�8D�"A߷ ��H��C-`����8�LRB� p��t���-8`��8�8Մ3� p��t���-8`ٴ�MA����7 �� 1�$Ʌ R��A�RA Ʌ	X�T5V�C_!@ȗT(� 5�TB���4V`� p�Tr'Ҁ��΃	�S@�R���N�8S�`1��8�n� 	ԃ� @ЅtŔC��`O SR% ���s�N �	��9P�``�B3R0���@�X�	5�`1�U� 5�N ɇ	ԃ��T"(Ү��wD0P�RP`N(A�@Ip ��Wq	ԃ	��@ߗR���N� �C�M%���D@��`2� @N$ �Q�> �����0��,8�`�M��1( ��8@ߧ�$�OCX�1��@N�1 N8�(`�c@���tR � �\,�� 1	�3M���N%% ���u R��A�RA �S���C@ߗϔNE%��	�8�`����?��u�H��0N�8�`	�8M�P�J����?��p�N2EX�	1�8M�`��P(`��8 ���sT	���D@R�   b)�w$��
(᠐�(�?������)k F��!.(/�!�&���a4>X��8+�`&� ��?࠮&_&&$'&'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[�   �  � �J�"~���� .ZY�X"�`&-J.
W�!#�(V0�v��?��U�""&+�J.�/�]� T�$^)�&�v�,.$T�!_bU`�!�S�/R!��~!!&��!bq*⠽�_!&*&$^)$t!�JQ7U�rP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!!.�Z�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��F.����&��� �択'8� ��/�����t����F.��� ����C	���MN �̀3`��R1`6N O�3�TN� PT0B# � �U� @��A5: ���D�E3: ���@	DA�0��0,�� � @` ��8�G5 � � @�N�� 5�N ��`1��	�8N�S�8T�           S	PRQ�	� 0CN���MM���ϋ���8��4� @��GLN� V�σN�`�a�4ԃՃ� 0Ń��C XQS %�D�΃T�# ��T5���8A	�	8�R2C � ��A3�8N`!�R1�� �DM�P��HG1L*�����DNa��C �D�U �#	�S ��A3�8�8��1�ϋ���8�NB�C�L �Ʌ R� 5L� Q�$ �D��U �#� 0�D�C��3�O��8DVC@��5DC�TɅR��C��R�� 8�(�� ��TO�#i  DT � � 0�� �   �P����� D8 0� 	��@	 D B �AD0RD  �P T�P �σD� �$ 0��@  P�  �����������������ҕR0@�a�A� @A�4 P � CA@6��# � 0U�� @�DM���C�P��C�BSR �BR1  y ������������TՀCO�3SQ �SF�N�Ƀ�ʆ��O��8J
��
.
���8@������/������O���&��0��&��HO��� �怀4ɀc�����&,�������������L� ����� � �ʀ&����x��h�����r

�����$ ���T���/����d����j��&�� 	�
���b�ؾ���   �� ����0 ���¬�b����d��6��D��ʐ���H����c ����4 ��D�△�P�䔒������     8������������)����)�������&�D.��b�����s ����2(���(/�ܢ��d�����J��d��*��h��������!������⮮c�����*   �� � L B    �@ �>��`�s�RS�(�!�s�b(���J!q���k�8�   � �W��C���{�����3D)��ʉp�3D)��ʉ'��a�������D9����ݢ�!|�ԫ�����d��6� � H �ۢ�݂��d͊���  �������J� ��w)  J
�
��(��H���                                                                                                                                                                                                