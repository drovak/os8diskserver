����   -	 	 . - 	 /8  -   /8   :      	 	  	?     	- 	,  	                                                                                                                                                                                                ��AT�0v&xş��C ���G �   �� �� ������E�?D0   �&���(ˁp�   ���8 �t�C ���0���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s�
��� �v���؇?����� ��)��)���b��������������.�i�����  ����� ����r�b
�b��y����T���
�~�b�f�� �� �
�&(?�	�6�&	�0!����J����D���� �� ?�!��� 
.

������ ���_��3�� �� 4[�C�������4��4�&�&���2���J�/��"�������)�������i����&�	&����b	�i��)�`������
&�	&	(?��	6(?��
'
'���
�r��i Z�&�	&����q�Z�/���k� ��i��bi ��Xp���� ���$��(�@"ރI8�EE�55
�����	&H?��6	�	H?�!��/�	�!⠊������)���/������&�	&	�?�	����		&H?�	�	7�	���)�x������������r��r�b�bt����b	�j�
�	(?�
�	6�&�H?�!��/����@��b���� �/�%���� �S	��($�2������IB���q>��/�����(��
t����������i��/����"�������񛍍����� 	  ���	  ����� ������/��� ��0����0H����	�� 	�z�	��T�F��{'�+��D. b ��p�Yb?� ��U �CJB����?��5�5۞6P cbȲ�H.����/�������/��J��.	�~F.	'���H.���H.bF�&	��*�	� ��bg�J� ��n&��c���&��c���!>h?���&&���H��� �67'��(?���H�s �=m)<�&���;� 3������	&
&
q>	0?����ھ�{&H?������D��tCt�J ��c�������6�C�����)����?������i�2��C����� �>����&�c���(�8���k 
.���(� ����雰 ���3��ބ5}�S� ���"��"��* ��&��  � ���D�J� ��
'�
'��K��(��(� � @���(��� ��ް��� ��(��� ��ʺԈ�+ ��"����+  �& . � .�����ī &!�ʀ�Ժ���� ����ދ ��������3��Ɋ� � ����� �?���� D�� �߀d��6��Cڀd�>܀d�H.�
n޲h��ʔ���(�����ۍm�F��&�ۂH!��@/�!���ރ-֕� �!�⠲�܅-�� �����-��"��҂��ʀ���K ������,��/���͏���K         � ����dB� !��(�?0B��!@�������}R�}�� � ����AT8A�ǁ�ǉ�E? ��sS`�CAF`&V`�BR1(-��Ƞ�5C"�@����A3DQ	��ON5.Q��wTL 	ϋ��� 0S��$�RA �3BR1 χ��T��WFճ�8D�0��GN� �Q�T@S��  �Rp��3�N��TO"� 3� ����!N.Q�Rq�	1�HF�`Sa�υu�uLD�����8�8VC@�R���>� ���N"S�`SRA��ԃń����DMS�"��w��3A5D(��5 �� N�@�S�"�Rp��3�L� �1��m�eT%�	3��D��EF.��Cp�TDT�C ���E��4��; �WFճ� 0�Wq� �D�0� H��3 ��A3 T�T "SRW�S�? X��s_ �sS`�TRmNB��� [NQT�'���T���  ����  ��  ''�'}������~ /�ӂ�*���
� �    <aR��b��&�K"F�H���&�P.��/�󩀀�����G���>��G+ԃ&�%L�G5S