����    � �   ? ?`��������  ;\�&��&v������C���["����&�&���Z�� @���/v�������&(/�&��,Z�9�?늬Z	��Y'����X����W�@?W���V��6U"�bT��'�c"�d�S���&�!.�?��@Z�W��!>��!��                                                                                                                                                                                                            ��                                        �� W                                    �!1@                  .墼��                  �5 �                                  �	Ł����� ��<����b�c(��	c(���	Ǒ�ʃ��*�<�� � Z	���  � � � � *��(ϫ �Z&�!�� > �   �j/�P�t
                        s��O/            ~�.�                               S���(� �8 >�&��&��i�(���������(���(/�@������i�����(/��������|�@��"��������"��&�*��b��������&��/� ���d�����/˃�~����n��b����j�H/��� �����/���}��i��� ���|˃�˃{�  3 �s��8����Å�q�����������K!�F��� �                                                                     �q�                  �%  M                              Ӽ� P                              [qp<���I ������ �,���,��7����A�K8������Ɂ�ȁ4ǂ�ɀ �4���Ɉ �9����P�� ���"��k            �1�                        ��#*#      ؗ J�                        � �                �� 鴇�                        �!V@            �  �                                                                                    ���      �e���                                                                                                                                                                                                                                          z��s                  e�0�G/                                                      N   �                                                 ��  �
      �� 4            es0 �                  
7�� ��<z&� "��D�!���� ��K�       �� �                   �� �  ��� � ����ށl�>���т���  �����  �����   �                        ���� @ �(����ЈЈ����� �        ��B�¨�Ӄ�� ����D��D��D ���b ���n��&����o��f�/��&�� ��b����&��0��&��3��@!�惃4��@��o��F���/��"J������݇�D �慢�/���� .��X���ƪ����V�������ݠ��������O�O���8�}���º�b��c�!��c����&��C��d��B���������������h��x��hb����t ����t8������      ���� � ��2 �����������"(���(/��������b���ޢĠn�Ħ��*��/���
V���r��f��&� ����s�����	��t�� ���0 ���¬�b����d��6��D������H����c ����4 ��D�△�P�䔒������      8  ������� ���)����)�������&�D.��b�����s ����2(���(/�ܢ��d�����J��d��*��h��������!��������b�����*   � (�����b�����(/����������&�JߔJ��&���(����/����/��Ӏd��"�����&$�(���(/���@�� ��˷�߸������*����� �����(��"�ނ����&� ����������L��� �&!��ޤހ߰����� � ����� �����}������������{���� ؅�� ��l�&��0��&��C��d��4������(��J�򹅄��P�H���8��4 ��D��خ� �   ��@���@/��"(��(���(��� /���@����o� � �� ����/��o�,��/�ʃ�˱����K��(�����(� .�� ���� �} 	 E ���8�           ��⑔j�8���| ����n�l��&��&��0��&��4�(��摑4��@���o��F�� ����J.��-��-���Dޠ�����"h����b ��X��J��V�������ݠ�����ު��O�O� � ���ȿ����'p�  � 8 ��}���v	P�nݏ_��F        ��B�¨�Ӄ�� ����D��D��D ���b ���n��&����o��f�/��&�� ��b����&��0��&��3��@!�惃4��@��o��F���/��"J������݇�D �慢�/���� .��X���ƪ����V�������ݠ��������O�O���8�}���~ �} �� �� ����6��C�����"����ݗ�� �� ����Ш� ��}���Ӡ��'�J>����/X��f>�������c�� �Ȓ���s
��Ԅ��/ԇ�����r��5�@/����c�����"A��`���'�㨆���  ���H����? 8�� ������&�����h ���7��D���   ��l��&؃����n��&�>�!��d��6��B��/�@?��4D�������
��Ç�؈��o��=�ꭀ�t ���� ��(����b��(��-�ꭀ������ԉ��؆������������ʢ�¨�������-����$�֚ pWgJ��(���o p} 8������j     �� ����&�挧��c��bD����b����d��6��CD�戃L���b��y���H�����ޅ��(/Ⅶ��B��&P�"���������Fޜ�(��Š/����� �� (�������F�����䪈PN��-����H/����d��JZw �{ ��ￆ�D��8 �/������������/�����b������@���ĸ�����-������8�?@�J�ֈ����ĸ�Ĉ����h����@�J�ɈĎ��ֈ� ���������� ����� � ���� !D���"��b �� ��f.��Ў� � ��(/����d��J\0  �  0��-��Ш���˖,��/@} ' }� ���f qi ga �.F�ⓠb� �(��q������E���   �� ����&��,��/�ʃ�� ���&��¯�b(����&��B��7�p��r�����q�� �          �	��쌇�

��s�F�H/�.��y��#��r��7�����7� �                   � (�������&��0H����&�>����C��d��6��L��&�����/ါ����H.�
n��h�����؍����m�F��&�H�a��-֫� �!��P ��鲅�҇���-�-��(��"(���k ����ۏ��촪خ����   � �     � Գ����� �       8����   P H  H H� � @�10(<H 2'?!	  ".2'?'  ,".
-2,,22'?!! 8".>2'=2"4242'?"   4".2'?*  9".2/<!   >
.;...I;?::<$ >4>A;''2 ??�B B <���������                                                                                                                                                                                                                Q8V��/�8�������m�(��@��|&8&8J.8����(���H/�J�V�8&��,� ���S��'�J>
��H.��J
��������u��(��!�瘨Ϩ �  � ���J^
�?H.��J
��� ��J.8��8�c8V�k              � g�P�@ ��� ��\�_"VU�2d� p �     �       �       �       �       �       �       �       �       �       �       �       �       �       �       �     띓��@��������Ӎ� ������?�!�}] c��   ��U�����D �B � ��                                                                                                                                   	 	                                                                                                                                                                                                                           � ��G��"����Z� �	�����  �	�Ԁ��	�� �� �� ��  (����/�ؾ���(����������  �   ��6��C�b�����2������    ��F���b���k �	�?����{�O�MN0 �3� 0��[               �T^���?�
G~T�����Z  ��������� ���|����� ������7��������&��2����Κ� ��㚣 ��U�� ��ۚ�ӳ�-�����-��� � S	Ut�DAN�!�R���DN(�A3� 0BT��QIu�NB�S�n �LS!ЃE:! �LS!L�TD� �                   �y�c�VG�V��?�������FN���&��,��|��C����������i�����i��������(������I �&���� �����,��|��K ���k �	󼳼�I���h�/��(�� (�����?�踩�h����b��x��b���暫�)�۪��+ ���<��K ���d��������D��� ���޴ � (����B���ǉ������˛���������� 5�����(���ɀ �5���K���< ����F��C�A�s �TEB3R �ϋR���DIV�8��4� �A q��@C1	�S                                                         �(�Ӏ��? ��)��7�����'��'��+ ���bg��J� ��]�R1��� 0���R���D�E���PL� �?�4R���D                                                                                                   ��:-^���������� � ���� �ᆢ��b�b��ǉ�Ȁ���<(����b��/��������"�������&�����* ������� ���ǉ����/��� ����  ����ӇD���&���ֈ������� ��� ���d�(?ֲ���J �	����$��+ �            � �����`�� xE���/�������2�����̨�� 7�����2(����/�����~��x����� ���ɀ ��� �� ���É����������'��'����:��̀`Sr�݀��0�H��A�3�N�G`����d� Љ��Y��A qO�3�T                            ��������%�V]y������,������ ���Ǹ��b�ψ������������� ���F.������&����&� .��&��"�Ղ�&��)���ւ�������փ����D���� ���&��(��J� ��р�� �       ���"��b�ڋ                � �@�?P	������S �U���	B  ���)��)����֞�����)�����)�����������	�����O~�Z<�? BYPG�                                                                                                                                       �  ��������� ���Ɂ�́����,���������#��ǂ�ɀ � �	��ɀ �6�	��Ɉ ��	���  ��	��Ɉ ��	��ˁ�É���ǲ��Ɂ ω��􃜁 ���ɀ �)�	���	 �0�	��Ɉ  4�	��������< ���� 4 ����� �   O��?�u �u8�� �G������&��&��tφJ����
�C � ��'��^��ǉ��8  ���� > ǂ��H� N ǜ� ���w��|���� �>����H �N�σ������Ɂ ΁��� ������&� �   ���(����s�����0�/��͉l����H�����@ u���� t
xG:� ��E��������������                                                                                                                                                                                                ��N�xş �
��������� � ����D   � � 4}���� F  ���&����p����d�ާ�و���������8����� �k�Z��O� 	��?�?PPS�������_K�λ��t*�F�	��	 �gP`v� v�s@�
܁�*� ��Ƈ`�D� Q�;�U���u������!>~�/�}�����������|y{z)yxrw��v�(��ui�9�{���ô��� �'��q��� ���ⲇ�{ࡨ��G��4�1�����,��7������
 t���4��c���c��͒��͛"���pb�l�.����& �� ����'8� ����/����tہ������ �0i͐��7g�����g�&o�ui'�v>�s7�eI�I�I��q�}��kL� Ө/�n�'��m�/�l��zY���&z9��|�wk&��Kkr|i{z)(?�z��{�z��jz)i"z|��=��f���Bf�e�F�&h(��d�(���@.c/����b����Ե�;�.&�����퀕�ba`��r�!�/�r�!�/�΢���r �!⠂�r�!⠂���/�r�������"��b��f΀h����V��&��&΀h�|�_D� 1^{��f��&��&���ċ ]	_��8Մ3 ^_Ο��4� 0^{_��L !� V^�����     � p� p ? ?`��؇��   ;\"��b�vi�/�����?��[�/���b��i�Z�� ���v���)�/��b(���b�Z�9����Z�	�Y�y���X侓��W�@W���/V��bU�&T)b��rc�&��JS�"��b!�����@>Z�/W�!��!.�?W��Ҡ���J��w ��p�dtZ^3Uf3u�����/R��^���/^R�����r�؈�_ӟS `^����'QP��u�C��T��F�� �� Q	Or� !�/Nr�!�/N��uS��T/�C/�  �M�R��e�r�U(`��/��L�r��s��_��� ^[�"b�kK !��hK��/�g��J�h��j_ğVC@^y� 3X�r)Xs�� ��QiJ��r�Is	u	S�T� �K !��hK���/�g�A�h��j��(��HZ�kv����(/�[��R�&&Q�b b�R�^�^J�r �riå���r��{�Z�	N�,G��Z���JyF�pE)�ρ �r��riH ��+ 6/"�"H.^ryL	��J��"�e���s�s)^���QP����MR�r���@.�/e���&Π/������D�zG�w��M���,�^{ �q�"��b�QiJu�C�� Ѓ RM^�s)^r��D�zG�wК�ۨ^ ���Á��� ��Cb��b�U�z����d�� �v����_ΟM@^0���"�b��a`��F�!!b!"⨔�|!�"�h�z)r����z)ք�rI �	r����z���r���||�_��  �)�)�z)�) �)#(/^T���&|_�υ` �^b�a`��r���r�Ȝ��ȊrI�	r����z֛]_��^�"�"։lց<$���;�SE)��ā���B)g퀸� ���	
�)_ȟNR�^b���s�$��c��{"�Б(?���������J��Ck���������⯆��6��C��d��� 6 ���_ٔ�RA�O���Abbg�J�R���bH/�!�w�/ۼ�"��bZ�����,�_�ω�ɀ���ZB)  ��B) 6 %�/E)� ˉ ��_����@^���%���ؑ�gvQP�uF�	 X PR��QO��&c"�b�F��ri�ZZ"�b�&!.�E)� Ɖ ��!.&�&����bT!��bc�&aʚ�F�a������r��s)�
c"ܶj!.ܠ/��!��&`ך��!��E����ܩ��!��&@y����&瘷(/^�����R�����?�����2�ET�����bfJi�_��� P^��~'?>'�='Z�'��~��~<%6��������j��JK T�Ӡ��bKt��������鵠���b��b�d�Ӫ��ŗ��;³ff�n��n��bhi(��b�@.��/���@.�/�u�R�� �_ӟNe ^k_ğ� @^��P?� ���E�����D�&�&����b	�b
�b�b�n"bia`��r��������/�F!�!""����rI���!!."�k��r�������!'�	�r�rib���.X�
'r����r�H 'r����r�J�s�������q:0J�(���ְ��fـfɔbF�t�����Ѽ���6d�"����+��^��y(/��&& &Or���r�Zs��`ryT	U(q�F�ri9 �+\�i�!���x��������'r����r�H �'�!���w���?���8r��{�(�e�(��7L)ri���r����V�j�������������� f�U�u
��_ZB) �6?2�5c?�&wB) �4E)��ʁt�4E)��ʁ��EB) �3Ų����B)o�#D.'�q�rU�&2E)�Á��E)��ρ���Z���&E)��É��� ����$�c�9���i�/9�"��x&!.��+T�v��'�F���i&�ir���s��������pE)� É ���7��Z���8ZsjY���m�K���l�����6�,���ˠޑ�Á�Z&�&@y���Z	��8������7��7��r��ǁ��#$���!.��wn�b �� �� /� /(��C�(���(/��(����R�)b�����J����#6�#+��B��z��(�2����"d!)b�\�[�&������@�� ��#�qG�/Q*@r��92;o��c&��@Z☀��C����!>��i@>Z�/����� ����c���b���?��B �?	1�( ���1�(��)�1�(7����?��B �?	� ��&��6��&X�B �?�B) ?ǛbryT	U(!�ri(/���!�:�&���8   � �_��� @^���7a��4�E�����p4E�����'�	a����.�cE��5�� 0�E�� �� ��b�b	c(���	cT/�(��µ&1B) `�J�	����à���M�9�e�� �����/R�#^k��/E)� �� �3B)  �1B) 6  .�E��'��$��ǁ_���D�L Y����@ ;��z���T駆���c��d��6��C��d��6��B�����É����D�����`��,��/��� �Ƒ���9��<�p�qK��?�_��TR`��HRC!? P9w)�v�G ��/������F���J�

�Ы���b����&,!�ʀ���԰@>��/��� �Nqs'�彠����E�S����Y� �E�x}� ��nc���J�?�������������)���������(����b�¨�����"�����Ĩ/���󀎰�8��4����� \��)��)ށ���{ �	!��܁<������D	�T5 ���Á���?�s8��h��)����$����)����f܊ � (i��� �q�? PU�� w�T��样⨟���&��"��b��l��6��É��ё,��t ��􏁬��&��"��b��l��6��É��с,��t��D����� d ��� �	��D����� ;��Ǥ��&��&��&���ߪ��&�0J
�
.
���󣚹��C���ȯ�������� �� �4x�������矣�����                                                                       ���                     ���� @ �(����ЈЈ����� �   �~	�"�*����� ��ӛ�T���;��<�	�م��� �  0 ���#            
7�� ��<z&� "��D�!���� ��K�       �� �                   �� �  ��� � ����ށl�>���т���  �����  �����   �                        ���� @ �(����ЈЈ����� �� �  �������⑔j�8���| ����n�l��&��&��0��&��4�(��摑4��@���o��F�� ����J.��-��-���Dޠ�����"h����b ��X��J��V�������ݠ�����ު��O�O� � ����   ������������� p ����� �"���� � "�*�����.�ZY�X"�`&-J.
W�!#�(V0�v��?��U�""&+�J.�/�]� T�$^)�&�v�,.$T�!_bU`�!�S�/R!��~!!&��!bq*⠽�_!&*&$^)$t!�JQ7U�rP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!!.�Z����w!�L���`���&!.(sV(�!�M�?���OP�a☞��`�PP7(V0(v�ZP�$!b!$�$$DP!�$0?K$��J�((m�O|�v �`&a'6�?��U����I`#�a�+ N�'����(?�"��&'O�����"2��~�t�##bp|��!�w��Vp.((#�JH �&��crG�/����� �P �T  ��.@V ~ ����C  R ��N��D�����N�p@����N��@����
��~�/ ����&�� �/��L!J�� z� �K�����5L�p@�� ��5L��@�� ��5L�q@�� ��5L��@�� ��5L�r@��  �5L��@��  �5L�s@��  �5L��@��  ���2��p�� �2��q�� �^p��
 �^q��
 ���� ����$� � ���� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 