����  �?/?7?;?=?>**************????              ?/?7?;?=?>???/?7?;?=?>**************b "/!>##/  "?##?#?#?"?#'!?  8!! ' $!! ' 8#?   0	! ' %!                                                                                                                                                                                                   �;`.:" � ���/�� �� �� �� �� ����D8�D��3]��- 7��h� xP�w�T�3�@  1��"�                                  )? Qe �� �� �� �   $ ����ݞ������������������� �����/�%`�,D�4�3�5�6�7�8� ��� ����� ���� ����� ���� ��ߥ�K ��� ��� ���� �߷�K ����T�Jl��������������P)���& ��J�Ā�O)�_�n �bD�.Hs�b �J��"�*n &��,� ��g�Bl���YB�A@f��@��A���'Y�BD&Ei��D�JE�JU����������������������&P�Ě ��ʚ ����"�i���� ��ޚ���/�-��b�p�   �
�@.b/�F�u��#��r��� 1"��#&O)�B�A`b@Ad�@�����ѕ������^������o� ��^� ���$&O)�B�A`b@Ad�@���̚������������&�� ���] ��_�bQF�u�7� �P(/i �Oy��m�L#� �JB �I�I]  ��I�^ ��I_  ��I�` �� �I�I]  ��I�^ ��I_  ��I�`(��� ��IIb] ��I^  ��I�_(��I`  ���� �I�I] (��I�^ ��I_  ��I�` ����69����B��X��JB6)b6���A&(?�6�����L�MgbB*b;;b<lb.dr��s�NrKhb:%k�K�MNbLgbB)b;;b<nb.dr��s�hr:%k�K�LNbMgbB+b;;b<mb.cr��s�hr:%k�C/�  �L�Q��e�s�S(`� ��̃�e@���?��b

�
���(� �e(�>�e>�ߋ ���������=�(�(�u� !��&��<⏄3g�B�nKMfL�oȐ�';&j.'b�*(;&k.'c�'��7h:&;<&<=&i9&��������YB�A@f��@��A���'Y�`�!�l �>���!..X.��h����- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0��3��� >`� ��B�CCd� �?>b!?�/�>!.=�?/9���=�JBD&Ei��D�JE�JU��_���� �l �l�������Y�:�����C�C�J<=&�%������d��6� � x �ۢ�݂��d͊���  �������J� ��w)  J
�
��(��H�� �}����s	�̾Ѝ�M������\�7��S")��ac=��X�%���Jx^_,��)R��n�C�r;٨�`sF_�4*��!��y�I�:$���b_z:Bі�(�~MD����jMr&�Ya�b{1��t�!yr)��B��vh:�)�~({ �i�`X`��M���]ٺн��H;�m���a/�s���C�L                                                                                                                                                                                                ����΃`�G��D�8 �U��1	ES�����`�LD!���D@R�8A�'����LD!��A��1	��T�>�_T` �GD�� 5�S`ǁ4`N2�TP?U U��� �LD!����΃`�GD�# �T? Pl�_R ���	�U��H��AM	�R1�D�����DD�� 5�A��@�H�`1�G���� ��@� X�@� X� � X�@K� X�@K��_��4��?� X�  ��_A�tBS��	�U��H��AM	�R1�D����� �D�8S�8��DDS�HS? ��N�A S�T��C�����E�UC�H�8��D�? @�o�D�TU�4׃���HST���S�T ��T� 5SA�,A��DR �T�o�p� � �1��m��^�lk�>nIR�>�n����>nI�� �� ��������޺�ފ��I�q���)����������K ����� .��d��J��d� �    C0 �� Hމ�R�. � �^��� ��߿�����}��i�P� PH���o  i�H�00HH��Z��� ���  ,?�S_����[��[J�ZP JP�JV� � ���H0D0H��E���U������r��{ ���"�n��"��b���# �@?�&2����+ �* p          on� ^`��a�_]��b�01 23 45 67 89 :; <= >?  ! "# $% &' () *+ ,- ./              	 
   01 23 45 67 89 :; <= >? �L�a`�Ca���'n1���3ai�3��_�����1�J�3��m��^�i��L�� � 0M,ذ����[h<[,@A BC DE FG H� JK LM NO  ! "# $% &' (� *+ ,- ./     �         � 
   @A BC DE FG H� JK LM NO � �֚��{ܚ� � �u�t� e�g}�e�  �                � @���v�}�s����g���  �  !�@     ��{���������������U��U��U��U��U��U��U����  �  !�@     ��{���������������U��U��U��U��U��U��U�!���`/�����)� �X              ��� ����%��� ������1��� ��0�?7���-��� �~��� �����������8GF'�$GF'�8� ` �I G'�%E�G'�)� ��� �~��` ����߈�߈�_��X 'V�'T�'V�'8�� �`� IG'%�EG�')������^��1�J�2��m��ث >�n� պ �� �����������ߺ�TRN�!  P�-��N�R� �� �� c��