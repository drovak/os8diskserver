��� m E-. 4#0>>30 ?0>7??$ t   ?>=<;>:.   ;&'988!= *
8< '9
*.
< '9	
	.  272	6> /5.#  '4? '3 2>(.+  +1>(/0
+>('/.5   .2	'4? +2&   /                                                                                                                                                                                                  ����B�l��&�� ����ہl��D���������@.�/�ozN

���&���� �  `����"��b�D��  ���&��&����������Д�c�J
��

��J��0��d��0�(/���� @�������c(���� �0 ��Z
�d�6F��K����f��P�S� ��&��&����(���  ����� ����y��L�����������خ���� ���l��?��(����&�F.�����bP�Ⱗ���̍ �   ����K ���?���������������ȟ��"����(/��튁�9� ȋL�W�  �9?P@��;PU� �:�P� �!�淸b��k � ��l��&��/����O����F.�බ7�J.
�����r��d��J��)��������d��'�O� �   � �   ���ŉl��0��&�?� ��,��/�˃�� ��/�ǲ�����г��&��+��S`Q	��  	a>�/�	�a�O� ��}����� K ��� ��������������9� �� �������@A����)����� ���&�'�&�&�'�j �	�/������c��c@�����z
�
����i���    �		���&������������&�à����������X.���O����PGU�`+fD�D]bH(��A]���
V:���g���'�y�&(?������̨/�������������� �	����'��0����>�����0�����?��� �������?����������)����i�ȿ��̄J   �i����"���'�J� �������t;�OYw�F5ُ��`�P� ��� ��W�������ȀF]ՀG��&�v���� �(/���(���&�"@������&���f��fрo'�B��/��������'��B����'��������'��)���&�'�J������'��)������c�/ߠ�&���z   �������`��������M�� [Og�r�ce�GM� Г&����&�(?�۹  ���I   �	���&�J� ��F���
��J���&�(?�϶��&��9  ��ȼ���"����X���"��w��#��y��w������	� ��������&�9� �����/�в�i���٫�����&]����ߙ�����ʆ���1�y��;uO�~       P�@�����  P                                                                 ������&(?���a��o���J�#��{� 0E�d ����ܣ���������/BD���������K�J�g��G�Y����������b�c(���s(����2��n&��?��C�~t�J�&�������� ( ��
>

������J� � �  ������ ��f��&��c(��@������dǀ��"(���(����J�ڊ��"��� ����)����� ��� j]��P?��I�O���ŏ����������&��b@����	cd6��(���c�c�c�cb �c(��!��a������    ������)� �� ����)�/�)��&�J�/������!��&� �����)P��_���ȚB ����� b��A8�.�(O�@�\d��	�������Ϛ(��Ǡ/����Ǣ(���&� �(/����(����������ǂ������ �@������&��)�������'���
.
���&`?�(���Ӏ��J�Ө���������� ��)������+����	H����v�T��    O�d��WO]�8;���`�Yt��g 
>

����� ��(���������H.� ��(/��(��H����)��������� (�����Y�F.���	��)�
.����������7� ���i
�   �������������  �   
��"�,8�HW�er��b� � F / A�8U��� �@ ����z
�? �8�`3���5TXL@!	�3σ΃�NL�_ R��A	5�8L@!N$ RQ��DL�_ �� �SNTT �Q 0���� 5`	��@�`6��  MATR`N �L�lL_! L�1 �0��4	��T [���p 	��@�`6�8VC_ 	���`Ra��D &!�ʀ���\���w��w��������c(���� ���J���c�h�bb��s�h��� �  ���� �  �����w��)젞��w� ��(?��!�� ���c���� ������'��'��� �a������;��D������O���C����c>����f���G?;��]d�K�����G��&������� �����6�	&	(?���&�	�b(��`��/���~��7!.�/�/��!�b!�b!��"�����S����2������grwr�u��(����렞�&�	�� �R`O`eՅD� �!.�/�〹݀��:��۔�����u��݄����r(/�������s���ؙ����H�����x���
  ��&��� �� Ж������������)��/������� �	���,��r��w��� �ϒD``k�	8�R1�DO�# m�R1��DN(-��	5�N2��σ`N2-�΃	�SN�!   ��� �����*� �·�Z�Yψ�Ov������i��&��&��&��&�?��Y�9  ���(��������?�����l� �   ���������&�(?֖�  �����  1���É�����	���j���  p ���"��b�盥�J����?�ʲ��b�j �	��ƴ]�� O�O�+c ��#��HƐ��� ��� �N���� �         �&��&��&��÷ ~��& ���J��쇁� ��MAA� ���'��0��'��'�c�l�� p���� ��/��5TX��C ��6��n��cJ
�
�� ����J��D�䢠����?���䔠�ꠄ��: 	7�J� �z�����?[���#H��ϑ������� y ��c�g��w��7� �����!>@/�
�� ?��
�J�
� /�	�
	&� ���É� ��� �������"��� ���c�����/ﵛ ��&��������Ɉ ��c�/Հ��/���k��dS�������	 ���{ �F8��;��oyO;a\���썓D��D3� ���&��'��0�����)�ӳ��P(q@�                        �72�                                                ��"�#                                                                      �	�Ф�