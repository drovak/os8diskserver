����  �@ �!;
2.   2:>29? *0
 8 2	*292	? + 
 $2.$        765/          
 *U5?/ > ? $2(  (< V ���������                                                                                                                                                                                                                                                   �	� ���� �޽Jݠ/ۅ�@������z
�
�⥂l� �  `�����&�� D��� ޓb��b��j��O�خ���˪��&��0J
�
.
��Ձ���<�����0��d��0�(/�����L�������<�����4ړ���d�X�'ӛ�t� \'e�'� � f��$ �	��  ���c��   �զ��������0�����0��z   ��b(��&�F.�����bP�Ⱇ����  
 ���K ���<��������/��)��������������!�����2(���(������ ���� )(�����:X"(������W��`����7W) �B?P@$��C$P��P��� ����F.����7�J.
�����r��d½J��)���� ��!.��b��b��k ���¾�l��?�������ā����<�����&��B��t���      ��0��&��;       ���*&[�& 
� `�6�' ��tׁ�� �/�i	a>�/�	�a���	a>�/��$ � � �$ �                                                                                                                                                                                                 	� �@ٔ�MA                                                                                           �            � ����dB� ��(�?��s��� �f � ������  � �� @� �"Ā� �? ���ѕ����效핈'��������
���� ����6� &��� b

�
���(� �(��� ���~"�(/��"���  )�"�����* &!�ʀ�� (,�b)�n+*f�(�*(B)@?Ӏ�)*B ��, / �� )�+��(�� )� �x�/�|��خ wb� �s߮!@� �   ���P�遼6����J&��ҹ~��~/}�-�H���� .� >����������r�J���Һ�}������~�-������ �   ���@�齼6��&� ���* ������o��"��b��o��&����&����!��H��J�r@`�q��
���-�-��aid��� 7;(��             ���b��6��&��ç����8��r��t��⢣d���� �         ��b����
.�দ&�� F&�� J
� .� ��n��i��/����d�ツ����&�I������&�J7J�6� �   ��� � F��J&Ja>�l�4�lv	��1	H�8�@< |{-�z&��~,ly&(?�����J��r��/�ɨ�ɸw�k��s��������e�Ѐ��q��!��v��}�� ��x��w�{�v{)�����!��� �u&�t�{ɛs&蠊�"����-${��-bc{���*-�J��* -���{-�{)�ɸzr|b{�(���ܠ���@ ���4H�������l�������"��"��" ��&��"H��D�J>�r���
��q0F�dF>p���*C
��CpD�d���C��D>� ��͛��F�����&� �!������&� � ���J��w"gw���   7 /W\�(7��� �=@�� �� ���4�����c�r@��3#63=N3W 0J
�
��o0�'���F���0����H.HH�c��t�n J
�c��
F�d�0����H.�dm0�'�N�J��n�F���D�0�D��dCl�
 ��D>��2�l���M�'� � /��xR()\()0a./�-�?8�������� �H��k@/�����i ������i   ��/��"��b�����/��&�!.������ ��k�&��&� �����O����H/�k�@����&���� � GJ
�n"""tGp J
����� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� W�@A�/ �B" G$ /�G�oG�"��l ��G�j�
ZDh�CpiCo������������lJ

�h�rF�gg7&�&� � �hgsg�&if0i�r"ie$(/����"�""G"GB""t���"GB�G�F�"��J$�/�G�HH�""7"GBqJ��$�/�G�F�"�:GD.""7"F�"�G�*����� ��&� ���D��D�%B���(/���&� � �eo0%dc

�
�ccF�&�!&���%%&$(/����!�!!C!j@��L�#�����!ⅅcH���!�!!D�!�

��o~�$����!r0F��!!CF�q��$����!>
��!n0F�!d!>�p�
!c!N���!!4��=� $ȉ��/�����b��i  ���) '�bb	�l	7	7	7"	c	s&r�y� �d� �����r'�n��r���b�bpJ
�irJ
�ghv�"&��� �	����&��&� �!�������H��k@/����j ���*Ձ,��K𠮁B†.c
�d0��3�@�^3̀/  (��
.r���&n ��&�D.�F.�b�p���"��bD��bF�D�⫪&M檀+    ��&K���&��/���"��j�b�H/��j�����"H����Fƀ���"���� )��)� )��"��"��c �� 9��C �� K������)� �   ���H�̭0ʰ �����@ ���� �(�b��r� �bp0���b6�&�&t�����r��r��~��y d���� bp �b�bb����� dऋ�亂�s�b��bk�he�2b�� �"(����/�ؾ�|�2�J&c�bbb�j!.�/�b�d����w����w�t������*x� x���� ��  %�l�����r�c(��c�lp (���~�  �����'�'m  p�Z
���r��b��i  `�e��p�dcF��b�d��� �����K �����#%D ��#&|E��#�b�#&##6#f��|��*C_�/��|i�b�c�� �k�h�P��$T�=A�d'D��]^D�M���<�&���'��ɉ���D$�c�#��0���b�?�������ھ����bcp �b��i d������s��퉜�&�?��bcp������ �o����� �ǋ�����*���~� ����bp0����䩈���雈�� �Pƀd��` ,E�$��=A�	楑����A ���������_��&��&��&b ?����~�@ `����b'bp0(�����~� ������y��� �l�6��(��p���� d��&�&t��߁n��i ���e��D����9�&����&�&�L&��(������恜� )� � �
�"d ��/%�������(����-��=��ƀd��@�� @�n��&�8l0�������������&��9�L����<������L�"L�e������J u t� ��   ��
.

������ �a �� ��&�&���
c!
���!>
�?��!
���"		c!
���	l0!
�����b��$���D�J� ������_�w��hߣ                                                                                                       �`A��� (P�p �����Prp�N� �P�ND!߃ �����C��wVC`��7��s��@V�C_! ��8q ���7Œt�8LTN�!���w�8�HL_! �TT �Q8�CR�� @�Nv VR�� @�Lr`� �QNQ   F.����&I���&�(?�Ƕ��0��7ƼJ    ������ܜ�̧�̬�̳����������
�I�KO�QG�IO�RT�aj�l ��k꠹��D��E�S����7RK�"�M)I� �(/���(���(/���������2(����(� �(���b�h����"@O��P��J�l .�|� ��"@�����P.�/��K ��b�nl0D ���2� ��'D���ᠮ# 0����#�##s�%&�%'�!.%�"�S���b��o �0�
F���W� �`� 89�n70f12f34f�6��&�ib(���(/���(���&�Ś����t�F���~b��/���0�/6�K34f��*7�K6�K0(/�8�19&���54bl46�K34f���&�"���#'���k�H+i ��@.��/��K�E	�g����k� �"@������%3�����F�0� `�b�lt����~�  :;f<=f>?f@AfBCf�z�c(����/�z�Eb.Fb/�i�"������(���H/��5F.5.5&�"���������/����&E.&F/&D&����D��i7�J.8&/9&8.&9/&CCB��/��(/�����z��j��(\T/���� ����-#�%� D� �/ 7�0����.8&/9&��&`&8�&9�&�~�
     �����������b�~�  ����������*45b��/5F.m���,0r1r2r3r4r�|� �P�� ���Z
�H� ���@�����i��� �
�~|i �/�]�)��!�t �G�/� �����_���K1 � �y  �� �ˇ� ��8b�9b��l~�    ���(�����)����:�!⨤�0�/��� d�:&�&�&�	&�<	�|�J��)����*��&0�/Ћ��~�0  ���"H��F�m��ǿ'��˿�j ��l�<HHb�� ��� ����������             x��� �0� LIU/�=� Cˇ� �(����� �F.��c���Hr�������r�����"��-�H������'��'��-���ȏ�~�-��?����t� ���߷��~�� ��~�-bھI�-������I���-��������/����������=����/�V�� �������   w����� @ }���� ���;  �� � ���&�����c�Jޘ���&��C�d��6��L�D��������&�����-��Р�������'�H���������"(���d�!.��&P���"���쀟����Fޡ�(���/����� �� (�������F������檀PN��-��N � � n� �t@��������D.8 �/����������&�������/��������P��젾�����-�������8�?@�J�J.����ǈ�ǈ�θ�Έ����h����@�J�J.����ӈΐ����� ���������� ����� � ���� !D���"��b �� �� .F��������� �  0       �
���ڠ����Ѝ�                                                                                                                                                                                                