����   @�
#,: -&: .<--<..,+#'?/      '62/3?}65 2-6/!5/ 4 ?/4=~ �B B (���������                                                                                                                                                                                                                                                                          	� �@ٔ�MA�':�!� b       A  �    � �� ���  +� @  �� @�   F
 I�    �`�     4   ����� S�O�^�UB��� R@� � ����dB� ��(�?��s�@: ��M��8m�e��a��$����?O����2���� ����������~��}����|���<�6�(?�{��&@>�/��������r��|��*�>�����}�����X~���)�}Á��F���~_����Љ�}�<�a�����'~�~�|z�<(��{�"�l�<�|���:���� 5�O� ��1 �0�/�/��Ԧ/��������'Z~�~�y��&����,  �ϣ����by �x	�� F����&��'�� �'��'�����r��ry ��y �)���r��s!��V����r��ry �)�	��y ���w�����耛 � �懃v�|���|���;�c��p�Q��l&!f#
o�h(�k&f f ��8,��> ��uɀ�4cJ
�
���8�J t (���(/�H���"���!�ʀu�� ��>�����7��0 ��s &����p !.s�/��� !��/�r���&�J����"F���b�h/��������&��"�c����r��'�'���|��z�� �6 .�t��l>�� ǁ���� 8 "�� ��@� ���&�����i	̒��
�����,�  ��J� ��� ���6��C��d�����������ہ �$ ���<����"�bqbc�c�t��� �������>���� ��b��r�}r�vB�L�Dp��&���r ���0����e�'��D^"��Z�#�� ���&�̚��/�ң��cςl� �  �Ր���b��"H����D�٢��&��D���׌*��������i��0J
���d��0F���оJ�����c����'��'��" ��ʄ&�ޢ�O� �   ��� )���, �����X�(������W��`����7W)V��7 /W\�(7���@U��7��� �±&ί�íJ��&ź��ͦ��ښH���&�?�
�

�����GùM�â ����2�����B��r��dˀ4�߀����&äJ� �ɹ&��J͎JÈj��ϟ,� ?Р`�     � ���-� �  ��ہ������-��ڀ��Ϫ���۠� �� Š  /��xR()\()0a./�/����$� 0�� �.�$ԃՃ�8��4� @N�$�CE�#҃`���@ R��C��S�� O�5�A��S MRMAN L#� ��C 1��P��p R�_P   ��2���|��z ��b�b�c�t�˫   ��Á�������) �ˀ� �� �� �� �� �� �� �� �� �� �� � ������f ���&�̚��/�ң��cςlԱ�  �Ր���b��"H����D�٢��&��D���׌*��������i��0J
���d��0F���оJ�����c����'��'��" ��ʄ&�ޢ�O� �   ����)����, �����X���?���Z������{ ������'����� �= ����\��#�ˌ�L�H>�������������&�㒠����2�����/��2�����7��/�����/��񀝁㢠����(�J>�����&��(�J��������(���j ��J>����������+鶟��� �#�T������� ��ݛ  �        �QϤO5��� ��#�f��C�1��6��\���M�=��   ��?���J�����H��������� ���d��4��?�����������k�  ��c��i��)�J>

�僳優 ��(�����������ր�(���������~����t� ������b��i�^�������a�́�+���:�܃��� ����R��Q��\��V����Q��࠰?��O�=� ��5�� ���i�ݦ���s��v��t��!������/��$��r��/�����/�������g��?����ɉ�ك �   ��&��d�(?���(���� F�����C����b�������b���q�ܯ�C��k�К�$��詌�   �����"̃������V�������Ѐ=�?�`=�#��\� ����U�fB��Lv��zL��j�:n�rD���&��%��)ή�r �(����(�����b������   ��� �&!̵��������� ���� ���?������ ��V���)� ���)��)� ��������ի�����±�ˠ�Ϡ�č����Рɠ�������"=͍  �ˣ��,���tO�3�T�R1E6 N E�LR@Q� 	�3����B �5 ��RA��D                                                                                                                � ��������������������������������� ��F����������&��?�����7���V5�Q�\��R$�������􃜣�����   ���������,��{ �	�������<�X��|����O��A��L0L� �CDD L�1 N2 E��  N � �$� 3XL`!�� p   D���Q�(�M��l#���⟽C��� � =� ������b��n��i�F>��Ϫ�0(����&��?�������t����!��/�.��7���f�� �	_����~��"��b����J��&��&���(������c��	(���/�������H>�����)�E��ݚ�����d��� �      ��t��J��CO ݇B�����#Qh�6	 ����� =̀�� ����i��)����£�b��b��h�#�������&���(�)������˿��p�������޼ �������g ���'�����7� ��ʬ�� ���&��C(���ƚ� ?���� ������c��d�����d��6ѠN��6�O��C���t���� �   ������ �@�ܟ��O�� ��=�                                                                                                                                                                                                