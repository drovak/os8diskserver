����  @ 2#*"**%
*; 2#2"*; 
%*20*.   ; > $8 !32-!8!<(*>

3		
<; <.*
3%3*3  	!! /     5,  >��������������������������                                                                                                                                                                                                 
 @ٔ�MA�� ���	    �#U(�" 0       Z[/����  � ��������������������7�7����������WX"�+� E� 3�8� � �
�? 	�  �@�  �%]I�    @�/��nsm&<�Y{ '�U��v���? ���?���R��` �H�j����&�̌(ϐ����(�,� �(���������)b��� (�����*�,� �(���������+b��� (�����,�,� �(���������-b��� (������.�,� �(������� ���&!l����(�����̀��(����/�, (�������� ��̀��(����0�, (������Ό(ϙ��1�� �(�����J��̀��(����2�, (������Ό(ϻ��3�� �(�����J��̀��(����4�, (���ƹ��Ό(����H�� �(�����J瀱c�%\�� �AP�CrR� 8         i� %"��l''O�%���&�J� b%�&�'�b!⠪��J�J�%���&�J/�����bbi %"��l#'�'�'OŹ����!�!b��fӒ%�&�%"�l ����!��/�����π���J�J� �  ����@�v��?�?`��؇��� ��!�!b��f��%�&�%"��l Γ ���!�⨡��H.
����������� � ���b%�& �� .����J �%�&��bt����*�!�(�5b6i %"�!b%�&�"'����� ��v��+��D. b ��l�Ub!�l!t=��!�z�<"�i;)�}��H/�(φ��>늤̜�́6� ���π��>�.! ⨠� /�>��J�KGK���>�6�� .����>ó�l'�>�%>'?%2??s�6d�>�  (��� k�[["��
 �A&B&@&	7b >c߁l�<	 t�ߢ�l�<C�|��&�<�|��&�<�|��&�<&�|�7�1�!�'&��'�|D''A&F& �����스�'�����(�i �&�%"� n f�� �J���9b �b	�b��l�<	 t�H� $b n t� �&�|!�&����J�J̀�O#�� �	 ?
� � ?� � ?� � ?������&!�@�W�W@���E��� 0�H>�$�!��� �����b�b�l�b��b%�&�!.�Hb�Hb��b%�&�!.��b��i �ށ< �"�!b�&!Ɂ��ä�ȿ����������� 0    �D� �������/�ߢ����¨���/ہ���˵�<��ˮ 0    � �
��(��&��J���   ����   J
�
��(��H��� ���6��C��d��6� B��b��b�b	�b��b%�&�Á	Ǧ�J��J���         �� %"��n�l����h�����%"��j��� �o'o .r�￾� �> ?��.���ʠ������Ӡ��������Ӡ������Ơ�����������������ɠ�������̠��������H��o$!$(/f�g�$@��!. b�&�����f���B%�&��� ��� 	� nt�	����	/�J��̤��& �&�I P�
J�!����!J� ��J%�"�Kd�H�K�k��N&&����M,��!M� �����!N� ������m����  X��������&&LLb����O�!L� ��JLP"LKd�H�K�k* P�$�!� �� �!�ʀ����P�&Z& ��,��_ ^_^6Ta'['X'T'/"�\b�k !^ / �!� ���̠�O�!�� �.���O���P�"��j(� �ɠ�������̠������������Š��������촄�&&ϊ���ϐ���ϖ��������ʄ��������������������������ʬ�ʄ����������ʬ����V(���������ׄ�؄������������堮��� �����ʀ�� ����������� �����V�� �����ʄ��V,����V� ��ʄ�����ʬ�ʄ����Ϧ������������������̷�������������� !��������V,����������P������  ���⬬䄬��� ��!����ʄ���ˀ�m������Ӯ��������ʬ�ʄ���ϊ���ʔ�ʄ�̴�������̛��������ʄ��(������
���������ϲ��Y� �  p                                                                                                         �U⇼l�̇ ������������X ���T�&������� �임������S�&�R"����������� !̳����V� ��� ��� �%�&!%"�dbebc n	�bI
J��I Jb"��|�<	ct���bb�l��O�ݢ%�&�%"��j��i�g��h�j���s������ ����!����ʄ�Ć�"������i r ����Y�ig'h��k&�̩�����W��Ķ���ٸŉ�ٸŠ������Ҡ������̠��Ġ������٠���������Í���Ķ���øŉ�øŠ������٠���������Í������ĸ�É��˸ŉ�˸Š���� ���f �&H�&H& �&����J���%�"��d�����&��ȃ�����%�&��D���ā�� �Ԅo$ !b��la!��(/�J��I J/�����%"��d� ��_'Xa'!R'�`'�S'� � 5 �3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�                                                                                                                                                                                                