����A   @�5-'  <;#':9;.6  0*?"-0.>  8000<(+'>+7< '>':/  2
$-: .': /<..<//-+$'?/      '62/4?}652-6/!5/ 4!?/4>~ �B B  ���������                                                                                                                                                                                                           ���v&xş��C ���       A  � � E�?D0   �&���(ˁp�   ���8 �t�C ���0���7�@ �� �� Zt1W����0 ?V������������� �K� 2��֩AR?�(�i�s���?�P�����/���� ����������~��}����|���<�6�(?�{��&@>�/��������r��|��*�>�����}�����X~���)�}Á��F���~_������zÁ�������"��s�/V~�~�|y�<(��{�"�l�<����V��O� ��� �0"�������b���������'Z~�~�y��&����,  �ϣ����bx �w	�� F����&��'�� �'��'�����r��rx ��x �)���r��s!��V����r��rx �)�	��x ���v�����耛 � �懃u�|���|���;|��僰�p�R��l&!f#o�h(�k&f f ��8,��> ��tɀ�4cJ
�
���8�J s (���(/�H���"���!�ʀt�� ��>�����0��s� �r� �l��' !r���� >!����q�"��d�����²F.����"h����/�����b�&��0��'��"�r�{�|�y;� ��cb �'��K?�ҁ����� �8"��!��@� ���&�����i	̒��
�����-�  ��J� ��� ���6��C��d�����������ہ �$ ���<����"�bpbc�c�t��� ����� ��>���� ��b��r�}r�vB�L�Dp��&���r ���0���쉼!�{�D^"��Z�#�� ���&�̚��/�ң��cςl� �  �Ր���b��"H����D�٢��&��D���׌*��������i��0J
���d��0F���оJ�����c����'��'��" ��ʄ&�ޢ�O� �   ��� )���- �����׳  ku�D)t&(?���H�s �=m)<�&���;�y�� 7:� �±&ί�íJ��&ź��ͦ��ښH���&�?�
�

�����GùM�â ����2�����B��r��dˀ4�߀����&äJ� �ɹ&��J͎JÈj��ϟ-�?Р`�     � ���-���ӱ�ρ����������݀���K���� �8)���|ly���a�S��*���{�x9��E���� �.�$ԃՃ�8��4� @N�$�CE�#M��`6��� �$��5��1� >O�3�T�� 5M$MNQ L�1 �4� 3���� �%_   ���/�|��y; �&��&7��J� � ���<������ ����ނ��d�����3���   ����   J
�� ������f ���&�̚��/�ң��cςlԹ�  �Ր���b��"H����D�٢��&��D���׌*��������i��0J
���d��0F���оJ�����c����'��'��" ��ʄ&�ޢ�O� �   ����)����- �����׳��?���Z������{ ������'��ڏ�> ����e��#�ˌ�L�H>�������������&�㒠����2�����/��2�����7��/�����/��񀝁㢠����(�J>���  �  �  �� �  ���(���j ��J>����������+붟��� �#�T������� ��ݛ!!�    � X�0�RϤP� �#�f��D�1��6��\���M�>��   ��?���J�����H��������� ���d��4��?�����������k   ��c��i��)�J>

�僳優 ��(�����������ր�(���������~����t� ������b��i�^�������a�́�+���;�܃��� ����R��Q��\��V����R��࠰?��P�>�!��6�� ���i�ݦ���s��v��t��!������/��$��r��/�����/�������g��?����ɉ�ك �   ��&��d�(?���(���� F�����C����b�������b���q�ܯ�C��k�К�$��詌�   �����"̃��@  b��� ���Ѐ>�?�`>�#��\� ����E�V�hBt�v��z�L�js�n��r�D���a�%��)����  �(/��������&��(��J� � ���� &!�ʀ������� �� ���c�����)� >�V��r��� �����Л ��� � ����-�����ց���0���� ��"���  �  �ˣ��-���tO�3�T�R1E6 N E�LR@Q� 	�3����B �5 ��RA��D                                                                                                                .25�9<�A �            DT � � 0��� ��F����������&��?�����7���V5�Q�\��R$�������􃜣�����   ���������,��{ �	�������<�X��|����O��A��L0L� �CDD L�1 N2 E��  N � �$� 3XL`!�� p   x����R�(�M��l#���⟽D��� � >� � ���l��&��&������F�옭��(�����cȳ���0�'��I��0!��������y�f�� ��_���7����&�/�夌���b�l�(?�����&��0�(��좠����?���H������E���֮��&�J��         P!݇B�����#Rh�6	 ����� >̀����� ����i� /�������&��&��&���$����(�'������*��փ������q�������� �����/�˵g� ���x�����{ ����� ���d�(?������ ���ě ���&ҭ6ҠN��6��C��d�����d���?��G��J�қ    �	����E/A�ܟ��P��!��>�                                                                                                                                                                                                