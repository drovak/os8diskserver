����  �= #!,-/48 "'+5	!+
!,0" , .!
!"""&"($$$$$$$$"$,$                                                                                                                                                                                                 � �i �8"`7�+    ��                 &!�"��� ~� � ���&&K� �      }�#����1� �9��zy�9�8 ��B��/��z�x�/BA�!�"�� #��W���`� �/K�"�
�F���� ����V����2�  H������ R>�����?�	� F�� ����bb �������ք����!⨚����Ȉ��J&�����&� �������oȢ�� !⨶����Ȣ��"(���o����/�&�����&�&��-�������Ш��������&Ŋ��� ���f�h���n �bD�.Hs�b �J��"�*_,$ �  �>� ������bwb��ߍ��ȅ�߄�ȅ��&����������ߨ�������n��ߩ��ȡ�߄�ȡ��&����������ߨ����&���� ���� �(/��� h��) ���	�(�) �������D�   ����� �(���� �� �����߀��� ZѴ A�qi^�S>�����b�m���������n�&�m���J�J���Ȁ��&��ل������m���������������������m������ȵ�������ȵ��&��ڀ�����������������mӀ�����������������S�(��RT)�!���s�g"�n�bQF�����Ū �� _!�|��&���� ������-�ߑ��������&������b�m���������m����������ߨ������������������m����ل������m�������&�������������������-�&��ڀ����������������M���*�JQ�*Y$�Q�M���+���tf�N9��_ !+�&��ڀ�����������������m������ȑ�������ȑ��&���� �� ހ�����Ƞ��߳���������n�&��ݹ��������J������������&�����&�&������������&��ڀ��J������������m�������:�� �`A�*��/� ��һ_��&�����Ȃ�������Ȃ���-�&����ք����� �������������m�������������������n��-��������/��������J����&��Р��������n��-����&�m����J�J������������&����� ���/Ծ�  �?� �l�@� �_o����b�m��-������� ���Ȁ��&�����ݗ�������������� ���Ȕ��&�����ݭ����������Ȫ���� ���������n��-�����Ш����-������� ����������6� � D �ۢ�݂��d͊���  ������k�?�g��� OM 6m!_�? ���&�����݅����������Ȃ���� �������������n��-�����Ш����-������� ���ȝ�&����-��������48f'+&�.�v0&18�u�#����A�/!..�/�.�0�J8t�.vb01hA/�!.��� .�.0d����.���//��cǛO@����ǜ� �` ���_� ?� h-�����"����������m�� ����$�����/���� �    ���-� � d��� ���-� � d����� ��
>

��(���H���(��0(���H/��"̈́� � ���&�.���b������J���   ��������� h̰��@����` ઺ ϰ0��@ � ��? �����������������ǈ��/������ ����(�� ������ �� &��� � �J� &��� � �J� &��� � �J��� ��� ���� �� �������� ���&���������R�&U&��K ���&� �(���z)�ﲠ��ᰰ �GIw�?����������������� �����b�m������b����ք���������Ȁ��&��-������b�����Ȝ��&���Ȭ���� �������&�����&�&����oȻ�� ���������b��������� �������&���� ���� 0T��T0C (��A�!��E������G � Ɲ@ �_ѫ������(��(��(��(��(��(��(��(��� ��r���b�bb򀞀��b� �����b� ���&�"ȝ��&�&�&�)����&�) ���)���&�) ��"b����������2(����z  ���=2��?Z@�(���:�
��9?�1#w w��f��f ���6��C��d��'�!>��?�����D���      ��c��d��t��J� �   ��c��d��篮D���    ���6��B��t��J� �U P ���6��B��b��c��t�O�Ҵ��J� �    ��RKm�_��"��b��� �@?�2����+ �*�{�=Ш�����o�n� ^`��a�_ � "� ���6��F��'� N��D���      ��c��d��b� ~��$��J���      ��c��d��'��D���   q ���c��d��'��D���    p ���� ����� ���� H̓TA@`ca���'n*���,ai�,��_�����*�J�,��m��^�i��   g�p � 0m,ذ���N�t�KG �,-&��#�����s��������������(/��������-䆱����!޸(/�!������-䆀��/������   ��s��t��7�.��y�������� ���7��C��r���8� ���=��Рr��g��e����� �� �� ��	������J̙�:�ed�8��?��@�9 � ��������������� ��� ���6��9�(��6��9 ������   ��� 0  ��)�(����� ���)�(�) �� ��) ��NTR � ��2 ���������) �����ٲ��� ��C�M%��� 0 ���C� �6:g >f
	   Z E��B�����Za� A�������) ������NTR��X��2 ���) �������C���C   ��������) ������	IS�8��C   ������q����� ���7��C�d��6�C�Ҕ�ë   � ��}�� >� pӛR!)O�JXO&^!)^!)R!)O�JQO&P!)Z^�!?��� 沞��`��H (� �,-&��"�����s��������������(/��������-䆱����!޸(/�!������-䆀��/������    ���6��C�d���������(������������ N����� >�F���������   �����%��� �� ����� ���y���?�	@  ���6��C��d��)�������(/�������Ǩ�ǈ�ǯ�� N��Jǯ���H����q�������      �������(/����������߿ �������� �������  ��b�!D����&�J.

���b�!D���� ��k e	ge�eY��}�_����eg�~e�=�� ٥Ә ���? 	D0��A� XGS�TR��CD�8A �MN ��A�RA��� 0NT"A	#�hS ��	 � 5�A��@MN0 ���R �C��$ ;�C Ĵ� KĄD�����A��D8D(�8R0��ăDD�ԃ�R��8R0D���HD(�8R0��ɇC8N`!�Gɂ NBԕD�O�N0 ��ɇC8N`!�G�Y�� E�8�L�Sh�$ ��3N�`�G��4� 5� E�8�Sԃɂ �D�3N�`�GR0D`�d� @ɇC8N`!�Gԃ�RD`���ɇC8N`!�Gԃ�RD`��C ��3N�`�G�8R0D`�d� @ɇC8N`!�Gԃ�RD`�ĄD ��3N�`�GR0D`�d� K��D ҳ��UDN`!�Gɂ NBԕD�O�N0 ��UD@N�`�GY0��D �S�`L@�SVɂ @UD@N�`�GT�8π3UD@N�`�G��4� 5� E�8`Sԃɂ UDDN`!�G�RD`���D UDN`!�Gԃ�RD`���UD@N�`�G�8R0D`�d 0UD@N�`�G�8R0D`�d� @UD@N�`�G�8R0D`�d� @UD@N�`�GR0D`�d� K��D ҳ��UDN`!�GՃ�R1	�/�A�8�8�D�`F�A� A	IS�8��Cɂ NBԕD�O�N0 ��	IS�8��C�Y�� E�8 L�Sh�$ 	I�3���8��4� 5� EN(A O1����DŃ��C �TP  	IS�8��C�RD`���D 	I�3���8�8R0D`�`�	I�3���8U��@ �S �T NR̓A�3G�S%�	EI�3���8�8R0D`�d 0	IS�8��CŃ��C �T NR��X�@1	IS�8��CŃ��C �PA��TR`�P�+ 4	IS�8��CԃT�`�ăD�,��D 0PX��4E ɃIU`�`C�SNR��R0R��%C���A�RA���TR@A�H��@G�S%��C �PA� �'ρ�A��H��@G�S%��C �PA� �'Ԅ��9A�4���GS�T� 5�A� A�'��E���ĕ�A��H��@G�S%��C �PA� �'��'��9V�A�4���GS�T� 5�A� A�'NTR0��'XNTR1��A�4���GS�T� 5�A� A�'NTR1��'XNTR0���L�C R��HS 	I�3���8T �8LC RQ��D�T@SX�`CNTR1 �׉��Y� 5�A� A�LC RQ��D׉�X��2�'5S� P�8�EÃ��# �TTS��`N5T0( �	�E��� �PA� ���X��2� 5��NQ҃��T �T`!҃��T �DT` ��R �D@T�`� ��� @��NQC��R  �T`!C��R  ���  \�C�D �H(�M�@P�-)��N���� �&!��"���� �=���(��Z�&;')��J�7�'v�&�,Q���K@����b��b��c��c����t��J�� �    1����� �� �� "/1����������������"	"
"!""$"(+"/1"7:"AH"NU"X["_�"��"��"��"��"��"��"��"��"��"��"�#33"%3'+35638=3@D3HS3TY3Z[3c�3��3��3��3��3��3��3��3��3�4DD D"'D+5D��D��D��D�EUHJUPRU��U��U��U��U��UԆW��w��w��w��w�.xJL����������"�, ���wLN��`�b���������������ę�ʙ����H�49 ;B DF ါ         ((�  pp�pp�pp�p(�$  >                                                                                                                                                                                                