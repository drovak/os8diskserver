����   � @    	 }:B K�����������������                                                                                                                                   �`C C� �W�R ��� 0�uN�T% �U3 Q ���VD �uN���@�uN�T% ��VD ��t�3C�8�1����C��G�G2 ȄF %�`C C� �WɇC8CcÀ1����D�4��sGN"L  ȄF %�UC5  ��@VD! �pݧ�W> nb����8� D�8�����3�m5���  0֭A�	��@�EE��� P�EE�	�  @�EE�D�T  ֔A��8 0֔A���F ֔A��PP֔A�����֔A���� 0֔A�	�1 L֔A��σD֔A��T֔A�C�	 D֔A���P 0֔A���֔A�B��A�|A��T�DK���M T��E����� �	�������������Iϰ���)��É��Ϟ������������ ����� .��d��J��d�j�      	�m� �D  ���� ����<Ȍ��Ū��É�� ������s� ������d��0(��@�
�

����(��@����)��J   � � � @�?E�C�  (�!" � ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    18}on�m{�| �>CGO]���y���۶��y�����g���ˀ��������d�򙀀�� � �	���� 1�mE��� P�EE����@�����Y@�EDC"��"��"��������6��H��h� �   ��)��9� ����������; �	�������)������ �	���/������,�<�����И��<�|��&�И��ÉF����ǉ���� !�/�����/�����/���������k    ��H �P���:�D   K����"��"CE"� ��(����`O   F��b��b��Ř�d���    ���(� .��bŧ����   ���A����������� ��� �	��I�Ÿ��b� �   ��b����&,!��"��ض-ڱ�Ҳ����    � �븀     � � J�~���#�;�~� �	 �����"ˊ �� ��� �l�Ao��n��&� �����?�����������)�����)�����)�Ò��)���ȱ�����ȟ�����y������E 8�LD  �� �C� Q�� 茀�TRN�!������ �� ���&��7� ������<���� �� ���� �	��� �	��� �	���� �    ������  �	������������ ���b��b��b� ���'��B���������&���� �!�澣c@������J!��!���"@�⣣K          �������TN"�  ���㉨���K �	 ��� ����� ����� ���ֺ��j�J���B����� �� � ���  �
� � �l�Ao��n��&� �����?�����������)�����)�����)�Ò��)���ȱ�����ȟ�����y������E 8�LD  �� �C� Q�� 茀�TRN�!������ �� ���&��7� ������<���� �� ���� �	��� �	��� �	���� �    ������ � �@ ��MA�� ���L �@  N����"L  ��WAN2�8D�R&B ���̚ ���$*�3��&��i���M������� u ?X�ڢ�* +�!���쪀 `    � � �� �               ���    ����M                        �W�2��vOfpwfx�bTYf_�i�/����:�~R�R� H
��&�	&	(?�z�z'�J��7��7��7��7��7�R yRb ���>y�H�R����&�"��>��L��/��b!����>��L��/���b��/�>��L����!"�#'�+ �(����o+�*�  �4���������_�?�S��Ey�}6-�3.�3�y�/�/�3�����Gz�+|�|� {{b!z⨢�{3)/�3�=��}6}�'�}{���� 5"V�"��"�-#��3,�3��3��4��3�F4��D��D��D��DO��Sb�����&��>�jw�x� ~���:R����nS�j@              - �A@ ���� ���"�:�w�Jx N�y��4�z�b( �3F�-�3F�.�3F�/�3E�4z��() 3�F��(+�{{b��/���z{b3E�4��(/�3F�-3�F.�3F�/3�F-�3F�.3�F��zzb� ި3�Fz�� ި3�Fz�� ި3�E4�4(��z6�&��&Ez�!��������3)E���$�4�?`����#����c�()�|�|P.@@�|�E|�({�z{b 3�F+�{�b|F�|/�zz!.{�/�{�3F�+{�{!.z�/�{�3E�|� ���4y��4�z�b((�+ �3F�/3�F/�3�F-�3F�-�3F�.3�F.�3�E4�M���b(0�  �3�Fy��4�(0�/3�F-�3F�.3�E4�=��!�z�<"�i;)_� @� M��(��l�0�  �p3iE4�M0��&��( �3�E4�y�/4M��()(/�  ��&�0�  ��0�p�/3E�4y�����&�0�2p��()(؞0p��3�F��(2�/�3F�-�3F�.�3F�z+i 3�E=���+��"�����b��k��"��b����!.�/�~������    ���P@� #��"�� E2�-��/��-�3�F.�3�F�����Gz�+|�|� {{b!z⨠�{3)Fz�|Bi���z{b3F�A4��()�P ����`&6���ba�h4�,��>-9þ��/��P�|.i3�F��P�zzb!�a /3E�� �������� �>�>	T��>����� 	A�� �
��)��&�@� �y �@� ���E.(��P����`6i�&�a&	&���+y	�z�a&�b&Qadb@N�P �P�a?�zz!.b�?���a|&b39E��P�!a���/�4���)�}��/4�4�=��׾�Ǿ���ݲ�!|�ԫ�����d��6� �   �ۢ�݂��d͊���  ��� � P��D���D���y>1� �@  P�g9P��|6|(){�j{,I-��/���{�/�Ůz{b3F�.3�F}���/�}���/�z&+|�|{&}�"����| {{b!z⨸�{3)FB���/���z{b3E��z&�4��|&�(�{o{|B,-���/Ϛ�{����z�{3)F.�3F�B����z&{3)E��z�i4 �?8 �M��8 ȿ�7@�35̢��`�k��~�`&�V�_&Z&9��X�b��{��H��4�H��4���4��1�����ǎ`�nVb_bZ9i�d�X���'�N����|9i�A95��4ž��"�`&�ô|�b(Қ+{�{!.z�/�{�3F�|-I��/Ӛ.�3E��ݴz�b(�z,)-��/��.�3�Eݛ@B   b���t�����f� L�H� �R(-�3�F/��+�{.i�{�3F�{� ��/���z{b3F�{� {{b���()-�3F�/��+{�.��{3)F{�������z&{3)F|��z{� |zb!|���{3)E���/��&��*�/�/��&��&6<�98�N?�k�J5֚4�        0/   /;: 	N@�?��� � 
`�  ��~Y��:~���}����V����&�@.HP��䑝��D.��+� � �{Od�.��~�~y���S��>��>ٽ�ޟt&Ht�G�}t&Ht�G
�H��G�H|�G�H{�G�Hz�G�Iw�x~	���G#�~�����D��S~i�:�Ol��5> +$>74+%.% 
>=>(+>0 ���/@ 6<�9���_r[lbk�/��_�kN@�k�J5��<9�8@�k�J5��4�~����?���

c(��}�/���qf�`����	&	!.�r&�r�s�b`F����b��icqbcq&c'	�J������"��*�3�̪�U�\�@�BA�C ��`� P�����cc&c'	�J� �    �	� .|���{�X�b@�����nV;i7���&Wi&Wj&�&)���-���,��jO�~����j��W�j�n`*��iO�~����i��_�[ZbY�jX�J�i����������&!.�/�>�L�G		Ϛ:���/��&~������>� ~	�:��O���i>ŝH��T&4 �               �A�Ei�^ �G�py�� �r��j�~V;iWd&7W�ehffgfWi&Wj&�*����\��i���~�����i�jV�/���Q(/��?�h�~�����්>	��>�>�~��:�Wi&eO�~����d�e�j�Ǌd�K�h�V�/���Q(/��?�_�[ZbYXd���`�~�c&c�2���� �                        ��f ���p����\��Wbj�bb�n)���Q��-i�0�+a�a�"��n`Jb���!a����(/g�Of~I�V���Q�/�g�������>	��>��⠿�>��>�>�&����n`�����>i->�3~�F����Q�/�>����bt&Jt�G��`�J�b?�tHt�G
�Ha�Q�K       �0-�`E{  �z��0�bL�j���~�����j�j�`�J��?��~�����Q�/�������>�8�㠩�>@��H��zQ�/�>�BJ�QG	�
Q(/��?�~��:��?�M����s̿d�M���6v�kLM�M�՚������ �            ��/   	��p@���  0lc,�P��2�1L��G��E{ ��w������(/��&�Pn�.��b:��(�(O���� .���F.�� �       ���/��K�� �kkb!l樱�_[&�` H
���&��&�Ƹ�ψ �$4�5ؘlk"����*_.�l�k�/���_�U�*���_b!_���_!.�/���                                 �	�8 lk"���kD.�k&k!.lb!�k�/���lk"����k�k!.l_b!��(�_�klk"����k�k�k����l�kH.�l�k�/�k�Ek�k!.l�j_!.�/�l�kH.!��_�k �� �����6M�� � �΀N�δ� �                                      �ƈ���� �X�f������V(/��O�Ǯ`���B ������"H�������"ǀn�Z&!.Z�/�Z�!����_D.�Zm&_�'�F>�Z��qr��3rrsr!>s�{   �����"F���
.��&��+��!                                                       {�z���� C� ����F��6��/�U��n��b@H�J��b��K����� ��!���6I �)��� � +
C+���c��F��4��ct�cu�b��f��&��&@t���&��u�&����t&�u&��J��/��� ��ڪ������"K����d��D��D�����"�v���`�����Ϝ�������� �   �H�� �C������‖6��"!��h��!���BK����� �
M����F��8��4��� ���� ��v�k�(/���@�K������j�¨��K��(��(��&�����b&��v�/�v��&��"���/�»�C��֣�KI�ݺ��4��b��n`����Hi�ݫ�v����� �JH�y ��
��@9��H��H �n�l��!��v�/�"��v�O�/�O��/i�p����0+��\}�"����P  J����`J�\ �� ��.���\����º>s�O�bD�� �    �Ol� �O�K�O�Ol�K�T����c.i c�� �                                             MҶ;@ ����6��Prn�c��/�����/���(/��.� +��]��2(/��.� +��^~�����S�J>ҝ������Q�/�����/�>��>ٽH�}G	�	�����/�>����Hn�G
���2�����2����>�JG�>	JG�>	J��H\�G�H]�G�� �                      �M��1 �
�� N�E0�H^�G�͉�Y�/�>���L[�G�LY�G#�͚���2���>�L�_G	(L	ZG	-H	`G	I	wx ��/�>� S~�����D����?�~����]��(/���(����/1~��:��M���2���� ����@	DA�0��0,�� � @` �� 5N���@1�N�� 5�N ��A����� �H��E+�P�P�-����P6�`���PP&P()��'��D�&�0��˚��P�n`��P"PPb(����rʁn0-��Z�,-��_�,��l�T&~����&�?o�JT�J����m�`\ P�
 ��\��j��E�4����b!�㚚&�	��R2C � ��A3�8N`!�R1�� �DM�P�ߦ���� �� @�@� �݀���ރ���&��*�ґ�b����&��ڑ�BT�ko�KT�K���������$p�p�-���*��/��.���Y��3��������,��s���� /�v�����v��������v���� ��v��C�߅tO�5A���	�P	�T  ��TO�#) DT � � 0�� �   ���9���E��o��t�0R�MT R�	��	1�8VC`�@�u�HRM TR� H�Rq�HT ��  � A��� 1�D �� 1��D�   �ńs���T ćVC`�HN�QT�  ߁q XN 1�dă`�`@�� H �R�  XS� T� @��c] NT" ��=8 	� ` R�$= �S� `_ ��E@ҷA- ���T� � �N  ���  �ST�`R��DT�`R��D �� @� � 1� �MuC��	� @� 0��sLD= ��@ͷS�$�8 A� @ՅsCa QR�ՅsCa Q�1L	�� �S�$�8��C���N�Rנ3R@$U�� W:���t�0R�MT R�	��	1�8VC`�@�u�HRM TR� H�Rq�HT ��  � A��� 1�D �� 1��D�   �ńs���T ćVC`�HN�QT�  ߁q XN 1�dă`�`@�� H �R�  XS� T� @��c] NT" ��=8 	� ` 