����  �C �  !< 
8!';
9?>(*%8';% : ';?7> 
 
';?6> : 54?3>(982?1> ;(8';;?';;?> 

0:?';	/? : .;/>(+ 

< 
>(-,+*/).y): )*3?<!>% > ! !??^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^���������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ m�
��D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �� �  �����}���v	P�n�_��Fn n�&J.
�����ȳ��������R.�i���b!�⨫�Ȁ����}�� %0����&W ��&�@�|"���J"��&���|����/�C��J��B(���}Ɉ � ���k   ��������������������������������HB�?������� �/ �� R�` VV�!�ڠ/�F����ڶ��r��x|b�i�(��m�������(��m(/�@��|��i�����m(/��������z�� �"�b� �F.��+�(/���H��bV�������m /���ڨ/��� ����� ��c�(�������F�� ���-�����?8��W��2d�pD�F�&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{ �(?��B6� � �gWq���� g�t��D����/���}�� $����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ���������  @��    �bH�
��bmF��B@���Pn�����彀�O��O��������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�׷�����2X��(?�
�

��������������o��R1��D��� N E��D� �@C� ����	��T P�ل�MA	O���� 0���/a� �&�	&�	��J�g�v ��V���T� � � �? ����  �&,
3��������������������������������������������������������������������������������                                                                                                  �����6��6���H }�� >Р�����c�c��{0(����bm�/mm"��bm�&��B�f��Ɉ }���k�c�� �������r`���O�֮��&���Γj � �w�?���&��&���?r��/�V��/����yN� PT0B# �텿��f����dw��DW�b��f�Dd#pD����&��) ���"�����)�J��� �	�����������{�
��*������/��"b��

d
(?��
1�����)
�9�������t�����������+�P���)�h� ���֣ � � ��  �/���/��?�˟�!��.�F$�@R��HH�V� �ɇ��`���o��W�>�����0�����S����0�����) ��������"������������y���E������B �A�B ��I��0�����������Ø�E��(?��c������9��`>�?�/������vÀ�� ��KW�x���P�O���Z x@1�Ywh�`��'����` 솀�����R��c(������ ��������+�����b���!�⠺��2�&�	&�&	7D�������7��� �� ��l)��  0��� ������ � ��@?ڀ��"�b!�@��d�É���Dܯ�����J��� ��=����c�/?�� �ɇhY����0�1������8� B�B��A�L���  0�L�	��@�L��� P�L�
�DC �vE�	�C0�vE�	�B1�vE� ����1 ��V���A �vE� � �	ct�᫣�z�����?[���#H��ϑ����Z����� 
 ��c�g��w��7� �����!>@/�
�� ?��
�J�
� /�	�
	&� ���É� ��� �������"��� ���c�����/ﵛ ��&��������Ɉ ��c�/Հ��/���k��dS�������	 ���{���F8��;��oyO;`\���썓D��D3̒�D3̒�D3�3�3�3�3�3�3�3�3�3�3�3�3�3��n��&��'��0�����)�ӳ��P(p ��b��&�J.����b�ۖ����J.P����U����"��b��&؉<�@.�/�����&��É�Ơ�� ��b���� ��ے�����)�����; �         �?����{ ����ů����� �KNUk�U������P��	�Ф� 8  ����� @3������ 0   !-6{|7z"7 �z�#�/g$�t� �u#    �� �      �}Ɉ 7	�7<��O�   � A�8� ����������������?���� ��!������ 3����� ���@� d�s���������������3-v �l�&�&���@~�����&7�㐋��	� ƫ ��  �����|�/�//D//D/�N�}Ɉ .�ؾ鐈!�l}�� ) ����|ɡ�b��hP��!��}�A /�
!�,ˀ�� BH��{�rz�~�y����z�xP�Փ���l��<� ���&�yÉ
Θ���}�   �
邼}I�  ����,�- /�w�|(_v*�w(��*�X�*ubtb"c!*⨡�"�J�/vs��"�rq)w|�p(�"(?o$��n�n�&!'&!,2���w�Po�m���hÂl}@���lt�$$bp ��X.��/!�x!����"k0�!'$�J'j;P"F�i�h�+Ii(g�**bf"&*e"!*bd(&!�;�ӛT�	݄ě���;��<� @������%!.cq9|&R!q�|o[  �%�&-bp(�b)�w$��
(᠐�(�?������)k F��!.(/�!�&���a4>X��8+�`&� ��?࠮&_&&$'&'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[�   ������i� �;`.    ������/� � .�� �� �� �� ����8����P���������� � U	UUUUUU!U#%U')U+-U/1U 0	5����G             � � #�49 I �	�����rM�i��^��mj�aE�LO�TW�Z]����0? ����E?�&�p����� �����s�nm�/��I�lp)�⾾d��m1�nm�2�q�lr)�⾾d�3�m4�sJ�lr)�⾾d�m�6���� ��R&#Q&%N&��&o�7m�8훀���brN�Ȁ�$N&K9�Q�J�Ț#Q&r)L:��R��������b� ��� ��f���<�ʁ�"�* ���� �������R&��&�*�R&��&�&�#�QbP�bO$bNoi;�m<��P�rN����$N&K=��Q����#Q&r)L>�POD���r)L>����$N&�x"!O�o�?m�@��Pr)N�J�$�NKiAO���P�N�&��&�P��!(?���ªd
 �  ��rL�B��R�J� �)2 ������� ���/���+&�,&���-�n-�-���-+D����+&�-��ڀⶱݟ,�����,&�-��ڀ��P_�����[�[m�Ń��C XQS %Z��}&Y&tā�X7�W2(��V(/�{�(��U�+T9��S(/�R�Tٚ! �s�g"�n�bQF�u�7� �P(/i �Oy��m�L# � ������Ҡn��b��bנnR$bNoiC�mD�׀�r)N�J�$�NKiER�����R&�ֲ��b׀nr)K����������բ��b׀nr)LF������&�R&�&" ��҃J��r��G����6���    #3  0" ��B�6I��&69����B��X��JB6)b6���A&(?����x ���)$N&�����/O&#Q&P&o�/m�0��Pr)N�J�$�NQd�����K1����#Q&K2�o�3m�5��r)L4����POD������� ��L�Q��e�s�S(`� ��̃�e@���?��b

�
���(� �e(�>�e>�ߋ ���������=�(�(�u� !���G� B � ���)$N&#Q&��&��&�����/�&�&�P&�O&o�/m�0P�r��NO�P�OO���߲�Ki1��$N&��&Q�J���#Q&��&��Pi�����O�j��&��&K2�o�3m�4�rL�5����D�����+3*H3* 0 �r���� 	A�� �
��)��&�@���E��G� B � ���)P&!�&!�&$N&#Q&o�/m�0P�r��N�J�$�NKi4���o�1�m2���rL�3���$�N�d����&�!�R$bN#bQoi=�m5�Pr)�N乀�$N&K6�Q�J���#Q&o�7m�8�rL�9��R�J������"�R!.�oi:�m;�r)�N��$N&K<����㹪    � ��t��G � o	��K��m����qs�pn�r��r)K��m����r�� ���)����i�!�Qb..bm����ݫQ����m)�r���J���   �������
&��&�!�QbmƚrQ�ƀ�
�6m)�r���J�۔������\ @ ����������������� ���&�yÉ
Θ���}�   �
����G� �� o	7���▔b�mi����J��J����P�� �   ��⪨b�mi����J��J������� �   �����b�oi� � ��  J��J� �  �   x����� ��H�������*bN�nQ�k��&$N&#Q&��K ���&� ������I��ŠTP P*e"!*bd(&!�;�ӛ�����ŀ�U�Ԫ�Kg   � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �����7�H.�S �"��c�U&U�"�����7��0J
�
���&�T6�� �X P    %%+d�%�] ?��� `!��k \��l)�� 0[� )�o(*f ��	6	 ?��������&�w  ����&��b

�
wभ�������� � �� P ��� �����"� �!��&!̱��� � ��(�("�� �&!���� "̲���!�*&$^)$t!�JQ7U�rP�~aa7(,2(OyN�a!�#&"�#�(�!�.!!.&�/�!�&�n*&M,6"%&!� @   �	�=���� �	�+�T�)�ז�0�S�)�ז���7Ub�����y����������K�j %e�H� 8 R���D��;  �0	�S �/�8�N`!NB�T�T 	�R1�D��� 0 �bc&�b&].^]&].^.^]b\���+                        ��fđW��e��U��� �	����������i���^�������������⻵b��b�i��b�V�DV�.�ix���������J� �� � W	�^��W�� ���f ���bH/�٤�ۢv�&�(/�v�F���׾k��*      
  ��`�e�Z�J��������T P           �   vĶU��X/)� �	������o�����o�����o������oǚ���o����inq��� �s˚o͚������o�������l �����o��������s�������������������������i�_���)�ז������D`R���C� ���V��U
	     u���ąme�]W���t m	�����+ �̉����Y � ���b����J.JJ�� �    ��� ��bFD�����+    Q����� ������b�mi��ǻJȹJ������� �   �������x���V��ʺ                                        � ��40���
7�Tp� ;� ENB�TXA��	�3��[�D@`�c ��HҠ3D��DT� ���H�`C�Ʌ.R �H��C	��R��KNT"A #A�3LS ��2 ��1HC�	�S1�X. �  ���� ��� ��������� ������%��� ������1��� ����<������ŀ�U �	�T���� ���&�����H�b�b	c	�t��� H��&� ��P��������|��������� �	�������R C��AG�8G,"S�T��CR� �	�Θ�ț�R C��AG�8G "F��@R�N�!�T1�C�. �QF�u�7� �P(/i �Oy�� �� ������U �	��������(��� ��� ��� ��������r��{ ���r��r�{ ��{ ���r��r��r�{ ���r�{ ��{ ���r��r�{ ���r��{ ���r��{�D��n�qǁ�ȶ�C�/�B�6I���%��T�$D
D��3õ3��3��3K93�=z 
  8 � K�	 �	����������ט��������������⑆j�C�S ��ԭԀKנK�m�`ô�`1�3�״��m`���AN NB m[Ӆ�l�pȄ18`��.8G�נK m�`�ŠT�D8S.   ����8�� ?��"�����'��J������ ��.��pݧ�W> nb���ߐ����U �$O&��(��'@/�(���&���m)�r�O�Jm����r�� �
������$$"�i�����$$"$N&����/m)�r��N䴏�   鐨����6쐠��#Q&���P�n$N&Pm)�r�N�JQO〮�P"PPb�H/���m�〮r)� � 5  ?� Q��PSɲNB� S9\8 �� �r)m������n��b�i�������bo��r�m��o���������������� �    �� �3;<���d���Z4�#�O��?�AE���d��ǁ>?A�E���dǓ�Z4�#�P����FiBښF�BޚC� �d���3Z�J������� ��w)  J
�
��( ��SRQ� ��*bO�b�nm9�r�O�Jm������� �� �� Ϯ �  ��  	���V��������ݳ�ݵ�ݷ ������&��&��&��&��&��&��&�����&� �����I �� �� �����K �� ���� �� ����                                     ����@� �� ��.&�^����i�� #�##bR�biȓ����$$"$$"$ .�Qfs�������Q�J��   � ����O�im��rO���� �m)�r����         �Q� ~��&�����R�K������ �                                               ��U��Q�ˆ�� ��&������#R&��&�ޜ��������"�Rd��� ��.��&�.�.��b����"�����︹"��/����+��    ��Ѡ�Ӣ��-i����-�����-��ڽ �|��N%�PE �S�  �0,�� � @` �� 5N���@1�N�� 5�N ��`?� ���׀���[ ��8���F��ⷮbF��⸀k   ��f��f��&͒��H?��������4��D�����k          �?d�
      �� ?�����t��J�����t��4ŀ�� ���&)�&��N%�	EI�3(�i 0`���  ���A� ����Ӡ  ��A� �`��Ӡ ���A� �� �0� �� �����������������'�������K ����� .��d��J��d� �    	C0 �� H �� ��/�� �������'��; ���6��C�(�@��

�
����0(���@/��"�۔� �   ����� ���&��'� �DT � � 0����@�?�	�� ��� � �� �����;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    ��}�tq�on�m{�| ����������� ���g�ܛ�ۖ��y��{��b�������d������� � � ��������� >��y����������J\ �7bޛ�@��
	�gh� f