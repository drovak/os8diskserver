����  �C �  !< 
8!';
9?>(*%8';% : ';?7> 
 
';?6> : 54?3>(982?1> ;(8';;?';;?> 

0:?';	/? : .;/>(+ 

< 
>(-,+*/).y): )*3?<!>% > ! !??^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^��^���������|�� G�,y�|Fn0��� ���i��&E0 i�Z
��c(O�|����d����Dc������� |�¨�����D�뢠����Ɉ ]�
��D����&��&��&�Ѫ�ߪ��&�0J
��
.
�������C��ȿ��� �� �  �����}���v	P�n�_��Fn n�&J.
�����ȳ��������R.�i���b!�⨫�Ȁ����}�� $0����&W ��&�@�|"���J"��&���|����/�C��J��B(���}Ɉ � ���k   ��������������������������������HB�?������� �/ �� R�` VV�!�ڠ/�F����ڶ��r��x|b�i�(��m�������(��m(/�@��|��i�����m(/��������z�� �"�b� �F.��+�(/���H��bV�������m /���ڨ/��� ����� ��c�(�������F�� ���-�����?8��W��2d�pD�F�&�`>E��� E��
���	&J&A�&��rE�/ @��f�����|�&�J��|�&O�������*���C 	�u�C !��H��	�r��J�&��d���(��!��F?0��0��7V F��'|�� /������"��s��{ �(?��B6� � �gWq���� g�t��D����/���}�� $����}���`�����c�Dc���բ��y�||�|	���t��J��<��r��z��/�m"�����'�����s�����'��'��'��D��J�� ���������  @��    �bH�
��bmF��B@���Pn�����彀�O��O��������� �v �  ��� ��0 ��� ��(� �&!̑��� �����c���J�׷�����2X��(?�
�

��������������o��R1��D��� N E��D� �@C� ����	��T P�ل�MA	O���� 0���/a� �&�	&�	��J�g�v ��V���T� � � �? ��e&<��KUgy�F����?��Dsp��d��8%W�Ȟb
�� �o�Ŀ����D�P��u�!�au���ٯl�M���o��0�yV��>뚒�����B���gz�O�0�͐�h�^�T����~u�m�7�ߗ�Fr�lPX-�9�l���m�Um���+~wW�<	����ԧ�����+                                                                                                                                                                                                ����&��) ���"�����)�J��� �	�����������{�
��*������/��"b��

d
(?��
1�����)
�9�������t�����������+�P���)�h� ���֣ � � ��  �/���/��?�˟�!��.�F$�@R��HH�V� �ɇ��`���o��W�>�����0�����S����0�����) ��������"������������y���E������B �A�B ��I��0�����������Ø�E��(?��c������9��`>�?�/������vÀ�� ��KW�x���P�O���Z x@1�Ywh�`��'����` 솀�����R��c(������ ��������+�����b���!�⠺��2�&�	&�&	7D�������7��� �� ��l)��  0��� ������ � ��@?ڀ��"�b!�@��d�É���Dܯ�����J��� ��=����c�/?�� �ɇhY����0�1������8� B�B��A�L���  0�L�	��@�L��� P�L�
�DC �vE�	�C0�vE�	�B1�vE� ����1 ��V���A �vE� � �	ct�᫣�z�����?[���#H��ϑ����Z����� 
 ��c�g��w��7� �����!>@/�
�� ?��
�J�
� /�	�
	&� ���É� ��� �������"��� ���c�����/ﵛ ��&��������Ɉ ��c�/Հ��/���k��dS�������	 ���{���F8��;��oyO;`\���썓D��D3̒�D3̒�D3�3�3�3�3�3�3�3�3�3�3�3�3�3��n��&��'��0�����)�ӳ��P(p ��b��&�J.����b�ۖ����J.P����U����"��b��&؉<�@.�/�����&��É�Ơ�� ��b���� ��ے�����)�����; �         �?����{ ����ů����� �KNUk�U������P��	�Ф� 8  ����� @3������ 0   !-6{|7z"7 �z�#�/g$�t� �u#    �� �      �}Ɉ 7	�7<��O�   � A�8� ����������������?���� ��!������ 3����� ���@� d�s���������������3-v �l�&�&���@~�����&7�㐋��	� ƫ ��  �����|�/�//D//D/�N�}Ɉ .�ؾ鐈!�l}�� ) ����|ɡ�b��hP��!��}�A /�
!�,ˀ�� BH��{�rz�~�y����z�xP�Փ���l��<� ���&�yÉ
Θ���}�   �
邼}I�  ����,�- /�w�|(_v*�w(��*�X�*ubtb"c!*⨡�"�J�/vs��"�rq)w|�p(�"(?o$��n�n�&!'&!,2���w�Po�m���hÂl}@���lt�$$bp ��X.��/!�x!����"k0�!'$�J'j;P"F�i�h�+Ii(g�**bf"&*e"!*bd(&!�;�ӛT�	݄ě���;��<� @������%!.cq9|&R!q�|o[  �%�&-bp(�b)�w$��
(᠐�(�?������)k F��!.(/�!�&���a4>X��8+�`&� ��?࠮&_&&$'&'^)!���'&D��(?�!�&�d�&���%2%+d�%�] ?��� `!��k \��l)�� 0[�   ����  i	 =�L��    � ��J$       �  �  !�@              ��� �������� ?  � �K��v�� � ���U��g��!~���� ���� �3?݇��!�� UU U(.U4:UBHUNTUZbUhnUtXQ XX(     � ����Qs��"��  @ �  � �������������=�Mk� ;�����&<��~�V(��%�� W!�~(/�%���
�:�<��}V)(��%�� W�!}�(��%�����:<��|�V(��%�� W!�|(/�%���
�:�<��{V)(��%ϐ W�!{�(��%ϐ�Ϫ:<��z�V(��%�� W!�z(/�%����:��캁�"�*n !I�D  g<��yQ)(��%� W�!y�(��%����:<��x�Q(��%� W!�x(/�%���:�<��wQ)(��%'� W�!w�(��%'����:<��Q�(��%:� W�!�(��%:�麪:<��Q�V�PW��(�%�L��:�<��Q��V�W��(��%[��۪:<��S� nS!�(/�%�j��:������"��<��Rv�d�T���%���T���%���P�T��%�����:<��R�RU���%��U��%���PU��%����:�<��Rv�d�T���%���W�H��%��ǳ�:<��R�RU���%ȑ�W�� �%����:�<��Rv�d�T���%ۑ��T�%ۑ�ۺ:�� ���?����C��m�L#�  $<��RR�U��%�,U��%����:<��R�T��RT��%��*�:�<��RR�T��U��RU��%��+�:�<��� &RiSS�SS�SS�SS�SS�SS�SS�SS�SS�SS�SS�SS�SS�U� N �J�� ��%/����:��6I��&69����B��X��JB6)b6���A&(?怢��<R�PR�U��%�����:<��R�T��ST��%���*�:�<R�T�����V)S!��(/�%���*�:�<R�T��S�!��(��%�����:<�RT��k��(̀��V)S!��(/�%���*�:�<��u&�&��۪%ϒ����:<��R�T�t&.V) �%���+P��:��߸�(�u� !� �?  �  �<��s&RR�T��U���.�V� �%��:P��:�<��r	&P��	6 .bV�QR�T��Wq� bp�/ "(��%�� � ����:<����PiR��T���%>����:������- !!�@,���h1�Zr��  ���?�+ ���Kr���� 	A�� �
��)��&�@���E��� 0��?<k�1������c��c�PiR �!Ti�P��&.V)R������=�L� Si����nQ�R�������=L�!�S�� !.!(/�H��*�@��%��ρ�:���k�����=�B���P�killb0V	lQ)RT��S��J�J lb�� �=L���J
� �d���3U���<e�fbPik��V)=G�k�qQ	�X) Z�Y��[��Z���&�JT����� �S!�k����!/=L� ��Z�P�V)�]�]�� & �JTƚ��� P�&�����܈�܈�$�$$�$5��ɨ������#�KZ�j����������?�_ƚ ��?��"�'���t#&#p)|�&����`�   ���6��C��d��6��C����!.��/��Ü�|��D��J� �    ���/�k������h�����)�)d(/�Ҩ�e���������k�����)"=L�k��О��b)&����K ��6�C��b

�
����(� � / (��-H/����� ��(�* ��'������ �ޠ �Yf�w X�=�L� Y�=�L� Z�=�L� [�=�L� \���=�L� ]���=�L� ^�=�L� _�=�L� Z�=�L� Y���=�L� X�=�L� ]�=�L� \�=�L� [�=�L� *���=�L� +�=�L� ,�=�L� -�=�L� .�=�L��/ � k	��k���$���8�/��)&)8&�*"��k�K�� �� � &9KZi����� ".�"��"��"��" 3=�3       k	��"�b�)"�k   �)"��c��dkȟ��� �	�����)���)�	��)�k���ˤ�/=L�����k �1��p�Y�f�JD�P �fh&��(gh&��(ce&��� �d(/�!�e�/�e��e&����K (?���0h'�5�;CUIOUU P[cUioUu P �  ��&(?���0e'����b�ctɶ�UU!U)/U      �+b�@n�.�����b�7���6�5ٛ   ��f��f��f�Yg�_3N&�/(f���*"&fPk��V	kQ�RT��S�"d�R�T��S�!.H/!(�)������� ����=iM�����v&k��V�QR�T��S�S�!.�/�ƪ���Ƭ���=�M��&�(�=�Gk����o �� &!��"��� ��(�ؠ�'�� �2����& 8���{�G��   ��   ���/�����"�=iG����k   ��� 4��g�g  � �	�v�ki�V	kq�  bQR�T��S��҂QW��J�S�b!⠻����� ��&��=�M�� �����"��
q���kU     	 
    �  ��/庼��@ ��'�m�k'l&B���a���f� P g ��<�3	&�2y���o�Pikl�l� V��lq 99bQR�T��S���?��	�|�J4��n&3	&��㠉�	�<if��㠉�	�<b!�jjb(����/�j���/���&�J�_�i�)�ޔ�����im=�M��i�Iyǚ ��n�b����B��� � 0	1�%�� ���Y�d� p� � �	<P�=L�k���  bX �Z��&�:�=L�k�llb ‎lq Qk�V�����&[Y����Z��R�T��Wq�. ��Q=�M��S`���_�b��/��^ʚa+���d�k���� X) Z�l�����lq Q�� �lq  ���D�l����&� �%�B�/%B���� H� �q�8�1� 5� ENQ�RD���PBI��4� p�	uI�3���8�1� 5� ENQ�RD���PBI��4� p�NuX�D	��R�H�R�A��wD�I� 1
XM��C��X߀�NqBG�S%��C T�R18�1�ށqLD!��Ņ�E	��R�HT "��߀ށqLD!��Ņ�E	��R�HT "	IS�8��C�߀ށqLD!��D0��A� P �d��X�8R0߀��w�LD�3D�8A L �N �3	��UI���EC�8�_1��w�LD��0P3X΅5�OB�N2�ɉDM_!��w�LD��4�C`��R1��C�E+��`K`ß��u��4�SɅEA��8UL@� p�Rq��C��4X�L@���`����� �O�3	�S�I��4� pޏsS`!N(L	UXAR�8D�F�Q��G�q�8�1�LDA �� 	���  ����T��A��wR���AGI A� ��	��0 `\�8U��D߀��p��LD!���A�A�8�1��w���LD��0A�R���AG� �D� I� 1XR0X���NB8T�$��wD�I� 1XR0΃_��Dp�HI �R��C� p�Dp�H OQ��LD!��� ER���AG� �	IS�8��C��� NR����7 �D�I� 1XR0΃`�G� ����LD��0A�F�����wF���� 5QA 51��߀�ޏs΃��TO�#	ESF����`1F��@N��8�#L���w���LD��0A�U 6�8��0`��W = � O� �P=  �PS``  PS�` �N �8�C2S��W�Dp��� ��R1�TU3P#�d	G��4C(-8D��C� p��t �T`�T�SN�  ��8�#	���-Nq ��8T�q[`�N�!`�N_
��wN �180 �ϖR���4��wN �8S��z���+�����na� �	�������������������������������� ����� .��d��J��d� �    
DC  �� H �	 �Ȍ��+ ������s� ������d��0(��@�
�

��ܓ�(��@����)��J   ���� ���&��'� ��b�����+Ϡ@ �?p?��=��!� � є�� ������;��A����b��c(����?�����J��?�����������K��C�����'��"��c��k    19}�to�nm�{|� g^@�IP�d����r��������i�����g���
�ܠ/����&��I������   � >��y�����������y���@��N������Q��@�?>=���݀�ݍ�������6��H��h� �   ��)��9��� ��?�>��� ��������ɔ������TRN�!   ���䲠����I�������̘�6��&�̘F.���d�� !�/�����/�����/��������������k   �`O `� HP���3>�  M����������=?��  F����&�� ��(�.�撆J� �   ��⿟� ����(��J��   �|�A�|��������� ���I� ������I�����b� �   ��b����&,!��"��ж-Ҳ����    ���&�����Ф�����f�f���� � 5R��TB � � 0����� �̸�����ʊЍ� � �� ��� �����A�����ɀh������������������)�����)�Ý��)�Ɲ��)����ȟ�����I�
�DC  ��LD!  ��N C�� �Q�> ����������� � 0U�� @�DM���C�P��C�BSR �BR1  y ������������TՀC� ��� �� �